`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Copyright: © 2019-2020, Chris Larsen
// Engineer:
//
// Create Date: 07/26/2019 07:19:00 PM
// Design Name:
// Module Name: fp_mul_tb_64
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module fp_mul_tb_64;
  parameter NEXP = 11;
  parameter NSIG = 52;
  reg [NEXP+NSIG:0] a, b;
  wire [NEXP+NSIG:0] p;
  `include "ieee-754-flags.v"
  wire [LAST_FLAG-1:0] flags;

  integer i, j, k, l, m, n;

  initial
  begin
    $monitor("p (%x %b) = a (%x) * b (%x)", p, flags, a, b);
  end

  initial
  begin
    $display("Test multiply circuit for binary%d:\n\n", NEXP+NSIG+1);

    // For these tests a is always a signalling NaN.
    $display("sNaN * {sNaN, qNaN, infinity, zero, subnormal, normal}:");
    #0  assign a = {1'b0, {NEXP{1'b1}}, 1'b0, ({NSIG-1{1'b0}} | 4'hA)};
        assign b = {1'b0, {NEXP{1'b1}}, 1'b0, ({NSIG-1{1'b0}} | 4'hB)};
    #10 assign b = {1'b0, {NEXP{1'b1}}, 1'b1, ({NSIG-1{1'b0}} | 4'hB)};
    #10 assign b = {1'b0, {NEXP{1'b1}}, {NSIG{1'b0}}};
    #10 assign b = {1'b0, {NEXP{1'b0}}, {NSIG{1'b0}}};
    #10 assign b = {1'b0, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hB)};
    #10 assign b = {1'b0, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hB)};

    // For these tests b is always a signalling NaN.
    #10 $display("\n{qNaN, infinity, zero, subnormal, normal} * sNaN:");
    #10 assign b = {1'b0, {NEXP{1'b1}}, 1'b0, ({NSIG-1{1'b0}} | 4'hB)};
        assign a = {1'b0, {NEXP{1'b1}}, 1'b1, ({NSIG-1{1'b0}} | 4'hA)};
    #10 assign a = {1'b0, {NEXP{1'b1}}, {NSIG{1'b0}}};
    #10 assign a = {1'b0, {NEXP{1'b0}}, {NSIG{1'b0}}};
    #10 assign a = {1'b0, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hA)};
    #10 assign a = {1'b0, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hA)};

    // For these tests a is always a quiet NaN.
    #10 $display("\nqNaN * {qNaN, infinity, zero, subnormal, normal}:");
    #10 assign a = {1'b0, {NEXP{1'b1}}, 1'b1, ({NSIG-1{1'b0}} | 4'hA)};
        assign b = {1'b0, {NEXP{1'b1}}, 1'b1, ({NSIG-1{1'b0}} | 4'hB)};
    #10 assign b = {1'b0, {NEXP{1'b1}}, {NSIG{1'b0}}};
    #10 assign b = {1'b0, {NEXP{1'b0}}, {NSIG{1'b0}}};
    #10 assign b = {1'b0, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hB)};
    #10 assign b = {1'b0, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hB)};

    // For these tests b is always a quiet NaN.
    #10 $display("\n{infinity, zero, subnormal, normal} * qNaN:");
    #10  assign b = {1'b0, {NEXP{1'b1}}, 1'b1, ({NSIG-1{1'b0}} | 4'hB)};
         assign a = {1'b0, {NEXP{1'b1}}, {NSIG{1'b0}}};
    #10  assign a = {1'b0, {NEXP{1'b0}}, {NSIG{1'b0}}};
    #10  assign a = {1'b0, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hA)};
    #10  assign a = {1'b0, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hA)};

// Broken code. See video for details.
//    for (i = 0; i < 2; i = i + 1)
//      for (j = 0; j < 2; j = j + 1)
//        begin
//         // For these tests a is always Infinity.
//          if (i == 0)
//            if (j == 0)
//              #10 $display("\n+infinity * {+infinity, +zero, +subnormal, +normal}:");
//            else
//              #10 $display("\n+infinity * {-infinity, -zero, -subnormal, -normal}:");
//          else
//            if (j == 0)
//              #10 $display("\n-infinity * {+infinity, +zero, +subnormal, +normal}:");
//            else
//              #10 $display("\n-infinity * {-infinity, -zero, -subnormal, -normal}:");
//          #10 assign a = {1'b0, {NEXP{1'b1}}, {NSIG{1'b0}}} | (i << NEXP+NSIG);
//              assign b = {1'b0, {NEXP{1'b1}}, {NSIG{1'b0}}} | (j << NEXP+NSIG);
//          #10 assign b = {1'b0, {NEXP{1'b0}}, {NSIG{1'b0}}} | (j << NEXP+NSIG);
//          #10 assign b = {1'b0, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hB)} | (j << NEXP+NSIG);
//          #10 assign b = {1'b0, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hB)} | (j << NEXP+NSIG);

//         // For these tests b is always Infinity.
//          if (i == 0)
//            if (j == 0)
//              #10 $display("\n{+zero, +subnormal, +normal} * +infinity:");
//            else
//              #10 $display("\n{+zero, +subnormal, +normal} * -infinity:");
//          else
//            if (j == 0)
//              #10 $display("\n{-zero, -subnormal, -normal} * +infinity:");
//            else
//              #10 $display("\n{-zero, -subnormal, -normal} * -infinity:");
//          #10 assign b = {1'b0, {NEXP{1'b1}}, {NSIG{1'b0}}} | (j << NEXP+NSIG);
//              assign a = {1'b0, {NEXP{1'b0}}, {NSIG{1'b0}}} | (i << NEXP+NSIG);
//          #10 assign a = {1'b0, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hA)} | (i << NEXP+NSIG);
//          #10 assign a = {1'b0, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hA)} | (i << NEXP+NSIG);
//    end

    #10 $display("\n+infinity * {+infinity, +zero, +subnormal, +normal}:");
    #10 assign a = {1'b0, {NEXP{1'b1}}, {NSIG{1'b0}}};
        assign b = {1'b0, {NEXP{1'b1}}, {NSIG{1'b0}}};
    #10 assign b = {1'b0, {NEXP{1'b0}}, {NSIG{1'b0}}};
    #10 assign b = {1'b0, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hB)};
    #10 assign b = {1'b0, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hB)};

    #10 $display("\n{+zero, +subnormal, +normal} * +infinity:");
    #10 assign b = {1'b0, {NEXP{1'b1}}, {NSIG{1'b0}}};
        assign a = {1'b0, {NEXP{1'b0}}, {NSIG{1'b0}}};
    #10 assign a = {1'b0, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hA)};
    #10 assign a = {1'b0, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hA)};

    #10 $display("\n+infinity * {-infinity, -zero, -subnormal, -normal}:");
    #10 assign a = {1'b0, {NEXP{1'b1}}, {NSIG{1'b0}}};
        assign b = {1'b1, {NEXP{1'b1}}, {NSIG{1'b0}}};
    #10 assign b = {1'b1, {NEXP{1'b0}}, {NSIG{1'b0}}};
    #10 assign b = {1'b1, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hB)};
    #10 assign b = {1'b1, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hB)};

    #10 $display("\n{+zero, +subnormal, +normal} * -infinity:");
    #10 assign b = {1'b1, {NEXP{1'b1}}, {NSIG{1'b0}}};
        assign a = {1'b0, {NEXP{1'b0}}, {NSIG{1'b0}}};
    #10 assign a = {1'b0, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hA)};
    #10 assign a = {1'b0, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hA)};

    #10 $display("\n-infinity * {+infinity, +zero, +subnormal, +normal}:");
    #10 assign a = {1'b1, {NEXP{1'b1}}, {NSIG{1'b0}}};
        assign b = {1'b0, {NEXP{1'b1}}, {NSIG{1'b0}}};
    #10 assign b = {1'b0, {NEXP{1'b0}}, {NSIG{1'b0}}};
    #10 assign b = {1'b0, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hB)};
    #10 assign b = {1'b0, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hB)};

    #10 $display("\n{-zero, -subnormal, -normal} * +infinity:");
    #10 assign b = {1'b0, {NEXP{1'b1}}, {NSIG{1'b0}}};
        assign a = {1'b1, {NEXP{1'b0}}, {NSIG{1'b0}}};
    #10 assign a = {1'b1, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hA)};
    #10 assign a = {1'b1, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hA)};

    #10 $display("\n-infinity * {-infinity, -zero, -subnormal, -normal}:");
    #10 assign a = {1'b1, {NEXP{1'b1}}, {NSIG{1'b0}}};
        assign b = {1'b1, {NEXP{1'b1}}, {NSIG{1'b0}}};
    #10 assign b = {1'b1, {NEXP{1'b0}}, {NSIG{1'b0}}};
    #10 assign b = {1'b1, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hB)};
    #10 assign b = {1'b1, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hB)};

    #10 $display("\n{-zero, -subnormal, -normal} * -infinity:");
    #10 assign b = {1'b1, {NEXP{1'b1}}, {NSIG{1'b0}}};
        assign a = {1'b1, {NEXP{1'b0}}, {NSIG{1'b0}}};
    #10 assign a = {1'b1, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hA)};
    #10 assign a = {1'b1, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hA)};

    #10 $display("\n+zero * {+zero, +subnormal, +normal}:");
    #10 assign a = {1'b0, {NEXP{1'b0}}, {NSIG{1'b0}}};
        assign b = {1'b0, {NEXP{1'b0}}, {NSIG{1'b0}}};
    #10 assign b = {1'b0, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hB)};
    #10 assign b = {1'b0, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hB)};

    #10 $display("\n{+subnormal, +normal} * +zero:");
    #10 assign b = {1'b0, {NEXP{1'b0}}, {NSIG{1'b0}}};
        assign a = {1'b0, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hA)};
    #10 assign a = {1'b0, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hA)};

    #10 $display("\n-zero * {+zero, +subnormal, +normal}:");
    #10 assign a = {1'b1, {NEXP{1'b0}}, {NSIG{1'b0}}};
        assign b = {1'b0, {NEXP{1'b0}}, {NSIG{1'b0}}};
    #10 assign b = {1'b0, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hB)};
    #10 assign b = {1'b0, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hB)};

    #10 $display("\n{-subnormal, -normal} * +zero:");
    #10 assign b = {1'b0, {NEXP{1'b0}}, {NSIG{1'b0}}};
        assign a = {1'b1, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hA)};
    #10 assign a = {1'b1, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hA)};

    #10 $display("\n+zero * {-zero, -subnormal, -normal}:");
    #10 assign a = {1'b0, {NEXP{1'b0}}, {NSIG{1'b0}}};
        assign b = {1'b1, {NEXP{1'b0}}, {NSIG{1'b0}}};
    #10 assign b = {1'b1, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hB)};
    #10 assign b = {1'b1, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hB)};

    #10 $display("\n{+subnormal, +normal} * -zero:");
    #10 assign b = {1'b1, {NEXP{1'b0}}, {NSIG{1'b0}}};
        assign a = {1'b0, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hA)};
    #10 assign a = {1'b0, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hA)};

    #10 $display("\n-zero * {-zero, -subnormal, -normal}:");
    #10 assign a = {1'b1, {NEXP{1'b0}}, {NSIG{1'b0}}};
        assign b = {1'b1, {NEXP{1'b0}}, {NSIG{1'b0}}};
    #10 assign b = {1'b1, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hB)};
    #10 assign b = {1'b1, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hB)};

    #10 $display("\n{-subnormal, -normal} * -zero:");
    #10 assign b = {1'b1, {NEXP{1'b0}}, {NSIG{1'b0}}};
        assign a = {1'b1, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hA)};
    #10 assign a = {1'b1, 1'b0, {NEXP-1{1'b1}}, ({NSIG{1'b0}} | 4'hA)};

    #10 $display("\n+subnormal * +subnormal:");
    #10 assign a = {1'b0, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hA)};
        assign b = {1'b0, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hB)};

    #10 $display("\n+subnormal * -subnormal:");
    #10 assign a = {1'b0, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hA)};
        assign b = {1'b1, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hB)};

    #10 $display("\n-subnormal * +subnormal:");
    #10 assign a = {1'b1, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hA)};
        assign b = {1'b0, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hB)};

    #10 $display("\n-subnormal * -subnormal:");
    #10 assign a = {1'b1, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hA)};
        assign b = {1'b1, {NEXP{1'b0}}, ({NSIG{1'b0}} | 4'hB)};

    #10 $display("\n1 * 2**1023:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7FE0000000000000;

    #10 $display("\n1 * 2**1022:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7FD0000000000000;

    #10 $display("\n1 * 2**1021:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7FC0000000000000;

    #10 $display("\n1 * 2**1020:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7FB0000000000000;

    #10 $display("\n1 * 2**1019:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7FA0000000000000;

    #10 $display("\n1 * 2**1018:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7F90000000000000;

    #10 $display("\n1 * 2**1017:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7F80000000000000;

    #10 $display("\n1 * 2**1016:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7F70000000000000;

    #10 $display("\n1 * 2**1015:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7F60000000000000;

    #10 $display("\n1 * 2**1014:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7F50000000000000;

    #10 $display("\n1 * 2**1013:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7F40000000000000;

    #10 $display("\n1 * 2**1012:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7F30000000000000;

    #10 $display("\n1 * 2**1011:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7F20000000000000;

    #10 $display("\n1 * 2**1010:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7F10000000000000;

    #10 $display("\n1 * 2**1009:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7F00000000000000;

    #10 $display("\n1 * 2**1008:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7EF0000000000000;

    #10 $display("\n1 * 2**1007:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7EE0000000000000;

    #10 $display("\n1 * 2**1006:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7ED0000000000000;

    #10 $display("\n1 * 2**1005:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7EC0000000000000;

    #10 $display("\n1 * 2**1004:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7EB0000000000000;

    #10 $display("\n1 * 2**1003:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7EA0000000000000;

    #10 $display("\n1 * 2**1002:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7E90000000000000;

    #10 $display("\n1 * 2**1001:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7E80000000000000;

    #10 $display("\n1 * 2**1000:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7E70000000000000;

    #10 $display("\n1 * 2**999:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7E60000000000000;

    #10 $display("\n1 * 2**998:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7E50000000000000;

    #10 $display("\n1 * 2**997:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7E40000000000000;

    #10 $display("\n1 * 2**996:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7E30000000000000;

    #10 $display("\n1 * 2**995:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7E20000000000000;

    #10 $display("\n1 * 2**994:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7E10000000000000;

    #10 $display("\n1 * 2**993:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7E00000000000000;

    #10 $display("\n1 * 2**992:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7DF0000000000000;

    #10 $display("\n1 * 2**991:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7DE0000000000000;

    #10 $display("\n1 * 2**990:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7DD0000000000000;

    #10 $display("\n1 * 2**989:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7DC0000000000000;

    #10 $display("\n1 * 2**988:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7DB0000000000000;

    #10 $display("\n1 * 2**987:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7DA0000000000000;

    #10 $display("\n1 * 2**986:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7D90000000000000;

    #10 $display("\n1 * 2**985:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7D80000000000000;

    #10 $display("\n1 * 2**984:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7D70000000000000;

    #10 $display("\n1 * 2**983:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7D60000000000000;

    #10 $display("\n1 * 2**982:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7D50000000000000;

    #10 $display("\n1 * 2**981:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7D40000000000000;

    #10 $display("\n1 * 2**980:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7D30000000000000;

    #10 $display("\n1 * 2**979:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7D20000000000000;

    #10 $display("\n1 * 2**978:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7D10000000000000;

    #10 $display("\n1 * 2**977:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7D00000000000000;

    #10 $display("\n1 * 2**976:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7CF0000000000000;

    #10 $display("\n1 * 2**975:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7CE0000000000000;

    #10 $display("\n1 * 2**974:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7CD0000000000000;

    #10 $display("\n1 * 2**973:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7CC0000000000000;

    #10 $display("\n1 * 2**972:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7CB0000000000000;

    #10 $display("\n1 * 2**971:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7CA0000000000000;

    #10 $display("\n1 * 2**970:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7C90000000000000;

    #10 $display("\n1 * 2**969:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7C80000000000000;

    #10 $display("\n1 * 2**968:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7C70000000000000;

    #10 $display("\n1 * 2**967:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7C60000000000000;

    #10 $display("\n1 * 2**966:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7C50000000000000;

    #10 $display("\n1 * 2**965:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7C40000000000000;

    #10 $display("\n1 * 2**964:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7C30000000000000;

    #10 $display("\n1 * 2**963:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7C20000000000000;

    #10 $display("\n1 * 2**962:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7C10000000000000;

    #10 $display("\n1 * 2**961:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7C00000000000000;

    #10 $display("\n1 * 2**960:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7BF0000000000000;

    #10 $display("\n1 * 2**959:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7BE0000000000000;

    #10 $display("\n1 * 2**958:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7BD0000000000000;

    #10 $display("\n1 * 2**957:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7BC0000000000000;

    #10 $display("\n1 * 2**956:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7BB0000000000000;

    #10 $display("\n1 * 2**955:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7BA0000000000000;

    #10 $display("\n1 * 2**954:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7B90000000000000;

    #10 $display("\n1 * 2**953:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7B80000000000000;

    #10 $display("\n1 * 2**952:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7B70000000000000;

    #10 $display("\n1 * 2**951:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7B60000000000000;

    #10 $display("\n1 * 2**950:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7B50000000000000;

    #10 $display("\n1 * 2**949:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7B40000000000000;

    #10 $display("\n1 * 2**948:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7B30000000000000;

    #10 $display("\n1 * 2**947:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7B20000000000000;

    #10 $display("\n1 * 2**946:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7B10000000000000;

    #10 $display("\n1 * 2**945:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7B00000000000000;

    #10 $display("\n1 * 2**944:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7AF0000000000000;

    #10 $display("\n1 * 2**943:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7AE0000000000000;

    #10 $display("\n1 * 2**942:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7AD0000000000000;

    #10 $display("\n1 * 2**941:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7AC0000000000000;

    #10 $display("\n1 * 2**940:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7AB0000000000000;

    #10 $display("\n1 * 2**939:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7AA0000000000000;

    #10 $display("\n1 * 2**938:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7A90000000000000;

    #10 $display("\n1 * 2**937:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7A80000000000000;

    #10 $display("\n1 * 2**936:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7A70000000000000;

    #10 $display("\n1 * 2**935:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7A60000000000000;

    #10 $display("\n1 * 2**934:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7A50000000000000;

    #10 $display("\n1 * 2**933:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7A40000000000000;

    #10 $display("\n1 * 2**932:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7A30000000000000;

    #10 $display("\n1 * 2**931:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7A20000000000000;

    #10 $display("\n1 * 2**930:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7A10000000000000;

    #10 $display("\n1 * 2**929:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7A00000000000000;

    #10 $display("\n1 * 2**928:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h79F0000000000000;

    #10 $display("\n1 * 2**927:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h79E0000000000000;

    #10 $display("\n1 * 2**926:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h79D0000000000000;

    #10 $display("\n1 * 2**925:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h79C0000000000000;

    #10 $display("\n1 * 2**924:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h79B0000000000000;

    #10 $display("\n1 * 2**923:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h79A0000000000000;

    #10 $display("\n1 * 2**922:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7990000000000000;

    #10 $display("\n1 * 2**921:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7980000000000000;

    #10 $display("\n1 * 2**920:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7970000000000000;

    #10 $display("\n1 * 2**919:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7960000000000000;

    #10 $display("\n1 * 2**918:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7950000000000000;

    #10 $display("\n1 * 2**917:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7940000000000000;

    #10 $display("\n1 * 2**916:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7930000000000000;

    #10 $display("\n1 * 2**915:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7920000000000000;

    #10 $display("\n1 * 2**914:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7910000000000000;

    #10 $display("\n1 * 2**913:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7900000000000000;

    #10 $display("\n1 * 2**912:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h78F0000000000000;

    #10 $display("\n1 * 2**911:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h78E0000000000000;

    #10 $display("\n1 * 2**910:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h78D0000000000000;

    #10 $display("\n1 * 2**909:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h78C0000000000000;

    #10 $display("\n1 * 2**908:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h78B0000000000000;

    #10 $display("\n1 * 2**907:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h78A0000000000000;

    #10 $display("\n1 * 2**906:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7890000000000000;

    #10 $display("\n1 * 2**905:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7880000000000000;

    #10 $display("\n1 * 2**904:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7870000000000000;

    #10 $display("\n1 * 2**903:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7860000000000000;

    #10 $display("\n1 * 2**902:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7850000000000000;

    #10 $display("\n1 * 2**901:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7840000000000000;

    #10 $display("\n1 * 2**900:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7830000000000000;

    #10 $display("\n1 * 2**899:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7820000000000000;

    #10 $display("\n1 * 2**898:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7810000000000000;

    #10 $display("\n1 * 2**897:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7800000000000000;

    #10 $display("\n1 * 2**896:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h77F0000000000000;

    #10 $display("\n1 * 2**895:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h77E0000000000000;

    #10 $display("\n1 * 2**894:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h77D0000000000000;

    #10 $display("\n1 * 2**893:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h77C0000000000000;

    #10 $display("\n1 * 2**892:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h77B0000000000000;

    #10 $display("\n1 * 2**891:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h77A0000000000000;

    #10 $display("\n1 * 2**890:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7790000000000000;

    #10 $display("\n1 * 2**889:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7780000000000000;

    #10 $display("\n1 * 2**888:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7770000000000000;

    #10 $display("\n1 * 2**887:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7760000000000000;

    #10 $display("\n1 * 2**886:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7750000000000000;

    #10 $display("\n1 * 2**885:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7740000000000000;

    #10 $display("\n1 * 2**884:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7730000000000000;

    #10 $display("\n1 * 2**883:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7720000000000000;

    #10 $display("\n1 * 2**882:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7710000000000000;

    #10 $display("\n1 * 2**881:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7700000000000000;

    #10 $display("\n1 * 2**880:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h76F0000000000000;

    #10 $display("\n1 * 2**879:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h76E0000000000000;

    #10 $display("\n1 * 2**878:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h76D0000000000000;

    #10 $display("\n1 * 2**877:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h76C0000000000000;

    #10 $display("\n1 * 2**876:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h76B0000000000000;

    #10 $display("\n1 * 2**875:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h76A0000000000000;

    #10 $display("\n1 * 2**874:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7690000000000000;

    #10 $display("\n1 * 2**873:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7680000000000000;

    #10 $display("\n1 * 2**872:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7670000000000000;

    #10 $display("\n1 * 2**871:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7660000000000000;

    #10 $display("\n1 * 2**870:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7650000000000000;

    #10 $display("\n1 * 2**869:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7640000000000000;

    #10 $display("\n1 * 2**868:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7630000000000000;

    #10 $display("\n1 * 2**867:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7620000000000000;

    #10 $display("\n1 * 2**866:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7610000000000000;

    #10 $display("\n1 * 2**865:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7600000000000000;

    #10 $display("\n1 * 2**864:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h75F0000000000000;

    #10 $display("\n1 * 2**863:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h75E0000000000000;

    #10 $display("\n1 * 2**862:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h75D0000000000000;

    #10 $display("\n1 * 2**861:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h75C0000000000000;

    #10 $display("\n1 * 2**860:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h75B0000000000000;

    #10 $display("\n1 * 2**859:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h75A0000000000000;

    #10 $display("\n1 * 2**858:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7590000000000000;

    #10 $display("\n1 * 2**857:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7580000000000000;

    #10 $display("\n1 * 2**856:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7570000000000000;

    #10 $display("\n1 * 2**855:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7560000000000000;

    #10 $display("\n1 * 2**854:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7550000000000000;

    #10 $display("\n1 * 2**853:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7540000000000000;

    #10 $display("\n1 * 2**852:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7530000000000000;

    #10 $display("\n1 * 2**851:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7520000000000000;

    #10 $display("\n1 * 2**850:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7510000000000000;

    #10 $display("\n1 * 2**849:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7500000000000000;

    #10 $display("\n1 * 2**848:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h74F0000000000000;

    #10 $display("\n1 * 2**847:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h74E0000000000000;

    #10 $display("\n1 * 2**846:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h74D0000000000000;

    #10 $display("\n1 * 2**845:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h74C0000000000000;

    #10 $display("\n1 * 2**844:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h74B0000000000000;

    #10 $display("\n1 * 2**843:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h74A0000000000000;

    #10 $display("\n1 * 2**842:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7490000000000000;

    #10 $display("\n1 * 2**841:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7480000000000000;

    #10 $display("\n1 * 2**840:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7470000000000000;

    #10 $display("\n1 * 2**839:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7460000000000000;

    #10 $display("\n1 * 2**838:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7450000000000000;

    #10 $display("\n1 * 2**837:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7440000000000000;

    #10 $display("\n1 * 2**836:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7430000000000000;

    #10 $display("\n1 * 2**835:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7420000000000000;

    #10 $display("\n1 * 2**834:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7410000000000000;

    #10 $display("\n1 * 2**833:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7400000000000000;

    #10 $display("\n1 * 2**832:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h73F0000000000000;

    #10 $display("\n1 * 2**831:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h73E0000000000000;

    #10 $display("\n1 * 2**830:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h73D0000000000000;

    #10 $display("\n1 * 2**829:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h73C0000000000000;

    #10 $display("\n1 * 2**828:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h73B0000000000000;

    #10 $display("\n1 * 2**827:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h73A0000000000000;

    #10 $display("\n1 * 2**826:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7390000000000000;

    #10 $display("\n1 * 2**825:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7380000000000000;

    #10 $display("\n1 * 2**824:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7370000000000000;

    #10 $display("\n1 * 2**823:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7360000000000000;

    #10 $display("\n1 * 2**822:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7350000000000000;

    #10 $display("\n1 * 2**821:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7340000000000000;

    #10 $display("\n1 * 2**820:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7330000000000000;

    #10 $display("\n1 * 2**819:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7320000000000000;

    #10 $display("\n1 * 2**818:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7310000000000000;

    #10 $display("\n1 * 2**817:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7300000000000000;

    #10 $display("\n1 * 2**816:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h72F0000000000000;

    #10 $display("\n1 * 2**815:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h72E0000000000000;

    #10 $display("\n1 * 2**814:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h72D0000000000000;

    #10 $display("\n1 * 2**813:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h72C0000000000000;

    #10 $display("\n1 * 2**812:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h72B0000000000000;

    #10 $display("\n1 * 2**811:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h72A0000000000000;

    #10 $display("\n1 * 2**810:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7290000000000000;

    #10 $display("\n1 * 2**809:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7280000000000000;

    #10 $display("\n1 * 2**808:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7270000000000000;

    #10 $display("\n1 * 2**807:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7260000000000000;

    #10 $display("\n1 * 2**806:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7250000000000000;

    #10 $display("\n1 * 2**805:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7240000000000000;

    #10 $display("\n1 * 2**804:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7230000000000000;

    #10 $display("\n1 * 2**803:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7220000000000000;

    #10 $display("\n1 * 2**802:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7210000000000000;

    #10 $display("\n1 * 2**801:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7200000000000000;

    #10 $display("\n1 * 2**800:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h71F0000000000000;

    #10 $display("\n1 * 2**799:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h71E0000000000000;

    #10 $display("\n1 * 2**798:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h71D0000000000000;

    #10 $display("\n1 * 2**797:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h71C0000000000000;

    #10 $display("\n1 * 2**796:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h71B0000000000000;

    #10 $display("\n1 * 2**795:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h71A0000000000000;

    #10 $display("\n1 * 2**794:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7190000000000000;

    #10 $display("\n1 * 2**793:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7180000000000000;

    #10 $display("\n1 * 2**792:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7170000000000000;

    #10 $display("\n1 * 2**791:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7160000000000000;

    #10 $display("\n1 * 2**790:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7150000000000000;

    #10 $display("\n1 * 2**789:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7140000000000000;

    #10 $display("\n1 * 2**788:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7130000000000000;

    #10 $display("\n1 * 2**787:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7120000000000000;

    #10 $display("\n1 * 2**786:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7110000000000000;

    #10 $display("\n1 * 2**785:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7100000000000000;

    #10 $display("\n1 * 2**784:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h70F0000000000000;

    #10 $display("\n1 * 2**783:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h70E0000000000000;

    #10 $display("\n1 * 2**782:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h70D0000000000000;

    #10 $display("\n1 * 2**781:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h70C0000000000000;

    #10 $display("\n1 * 2**780:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h70B0000000000000;

    #10 $display("\n1 * 2**779:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h70A0000000000000;

    #10 $display("\n1 * 2**778:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7090000000000000;

    #10 $display("\n1 * 2**777:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7080000000000000;

    #10 $display("\n1 * 2**776:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7070000000000000;

    #10 $display("\n1 * 2**775:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7060000000000000;

    #10 $display("\n1 * 2**774:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7050000000000000;

    #10 $display("\n1 * 2**773:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7040000000000000;

    #10 $display("\n1 * 2**772:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7030000000000000;

    #10 $display("\n1 * 2**771:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7020000000000000;

    #10 $display("\n1 * 2**770:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7010000000000000;

    #10 $display("\n1 * 2**769:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7000000000000000;

    #10 $display("\n1 * 2**768:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6FF0000000000000;

    #10 $display("\n1 * 2**767:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6FE0000000000000;

    #10 $display("\n1 * 2**766:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6FD0000000000000;

    #10 $display("\n1 * 2**765:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6FC0000000000000;

    #10 $display("\n1 * 2**764:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6FB0000000000000;

    #10 $display("\n1 * 2**763:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6FA0000000000000;

    #10 $display("\n1 * 2**762:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6F90000000000000;

    #10 $display("\n1 * 2**761:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6F80000000000000;

    #10 $display("\n1 * 2**760:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6F70000000000000;

    #10 $display("\n1 * 2**759:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6F60000000000000;

    #10 $display("\n1 * 2**758:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6F50000000000000;

    #10 $display("\n1 * 2**757:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6F40000000000000;

    #10 $display("\n1 * 2**756:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6F30000000000000;

    #10 $display("\n1 * 2**755:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6F20000000000000;

    #10 $display("\n1 * 2**754:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6F10000000000000;

    #10 $display("\n1 * 2**753:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6F00000000000000;

    #10 $display("\n1 * 2**752:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6EF0000000000000;

    #10 $display("\n1 * 2**751:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6EE0000000000000;

    #10 $display("\n1 * 2**750:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6ED0000000000000;

    #10 $display("\n1 * 2**749:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6EC0000000000000;

    #10 $display("\n1 * 2**748:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6EB0000000000000;

    #10 $display("\n1 * 2**747:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6EA0000000000000;

    #10 $display("\n1 * 2**746:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6E90000000000000;

    #10 $display("\n1 * 2**745:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6E80000000000000;

    #10 $display("\n1 * 2**744:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6E70000000000000;

    #10 $display("\n1 * 2**743:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6E60000000000000;

    #10 $display("\n1 * 2**742:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6E50000000000000;

    #10 $display("\n1 * 2**741:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6E40000000000000;

    #10 $display("\n1 * 2**740:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6E30000000000000;

    #10 $display("\n1 * 2**739:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6E20000000000000;

    #10 $display("\n1 * 2**738:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6E10000000000000;

    #10 $display("\n1 * 2**737:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6E00000000000000;

    #10 $display("\n1 * 2**736:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6DF0000000000000;

    #10 $display("\n1 * 2**735:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6DE0000000000000;

    #10 $display("\n1 * 2**734:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6DD0000000000000;

    #10 $display("\n1 * 2**733:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6DC0000000000000;

    #10 $display("\n1 * 2**732:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6DB0000000000000;

    #10 $display("\n1 * 2**731:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6DA0000000000000;

    #10 $display("\n1 * 2**730:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6D90000000000000;

    #10 $display("\n1 * 2**729:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6D80000000000000;

    #10 $display("\n1 * 2**728:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6D70000000000000;

    #10 $display("\n1 * 2**727:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6D60000000000000;

    #10 $display("\n1 * 2**726:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6D50000000000000;

    #10 $display("\n1 * 2**725:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6D40000000000000;

    #10 $display("\n1 * 2**724:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6D30000000000000;

    #10 $display("\n1 * 2**723:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6D20000000000000;

    #10 $display("\n1 * 2**722:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6D10000000000000;

    #10 $display("\n1 * 2**721:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6D00000000000000;

    #10 $display("\n1 * 2**720:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6CF0000000000000;

    #10 $display("\n1 * 2**719:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6CE0000000000000;

    #10 $display("\n1 * 2**718:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6CD0000000000000;

    #10 $display("\n1 * 2**717:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6CC0000000000000;

    #10 $display("\n1 * 2**716:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6CB0000000000000;

    #10 $display("\n1 * 2**715:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6CA0000000000000;

    #10 $display("\n1 * 2**714:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6C90000000000000;

    #10 $display("\n1 * 2**713:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6C80000000000000;

    #10 $display("\n1 * 2**712:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6C70000000000000;

    #10 $display("\n1 * 2**711:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6C60000000000000;

    #10 $display("\n1 * 2**710:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6C50000000000000;

    #10 $display("\n1 * 2**709:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6C40000000000000;

    #10 $display("\n1 * 2**708:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6C30000000000000;

    #10 $display("\n1 * 2**707:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6C20000000000000;

    #10 $display("\n1 * 2**706:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6C10000000000000;

    #10 $display("\n1 * 2**705:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6C00000000000000;

    #10 $display("\n1 * 2**704:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6BF0000000000000;

    #10 $display("\n1 * 2**703:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6BE0000000000000;

    #10 $display("\n1 * 2**702:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6BD0000000000000;

    #10 $display("\n1 * 2**701:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6BC0000000000000;

    #10 $display("\n1 * 2**700:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6BB0000000000000;

    #10 $display("\n1 * 2**699:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6BA0000000000000;

    #10 $display("\n1 * 2**698:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6B90000000000000;

    #10 $display("\n1 * 2**697:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6B80000000000000;

    #10 $display("\n1 * 2**696:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6B70000000000000;

    #10 $display("\n1 * 2**695:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6B60000000000000;

    #10 $display("\n1 * 2**694:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6B50000000000000;

    #10 $display("\n1 * 2**693:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6B40000000000000;

    #10 $display("\n1 * 2**692:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6B30000000000000;

    #10 $display("\n1 * 2**691:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6B20000000000000;

    #10 $display("\n1 * 2**690:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6B10000000000000;

    #10 $display("\n1 * 2**689:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6B00000000000000;

    #10 $display("\n1 * 2**688:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6AF0000000000000;

    #10 $display("\n1 * 2**687:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6AE0000000000000;

    #10 $display("\n1 * 2**686:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6AD0000000000000;

    #10 $display("\n1 * 2**685:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6AC0000000000000;

    #10 $display("\n1 * 2**684:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6AB0000000000000;

    #10 $display("\n1 * 2**683:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6AA0000000000000;

    #10 $display("\n1 * 2**682:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6A90000000000000;

    #10 $display("\n1 * 2**681:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6A80000000000000;

    #10 $display("\n1 * 2**680:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6A70000000000000;

    #10 $display("\n1 * 2**679:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6A60000000000000;

    #10 $display("\n1 * 2**678:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6A50000000000000;

    #10 $display("\n1 * 2**677:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6A40000000000000;

    #10 $display("\n1 * 2**676:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6A30000000000000;

    #10 $display("\n1 * 2**675:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6A20000000000000;

    #10 $display("\n1 * 2**674:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6A10000000000000;

    #10 $display("\n1 * 2**673:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6A00000000000000;

    #10 $display("\n1 * 2**672:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h69F0000000000000;

    #10 $display("\n1 * 2**671:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h69E0000000000000;

    #10 $display("\n1 * 2**670:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h69D0000000000000;

    #10 $display("\n1 * 2**669:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h69C0000000000000;

    #10 $display("\n1 * 2**668:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h69B0000000000000;

    #10 $display("\n1 * 2**667:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h69A0000000000000;

    #10 $display("\n1 * 2**666:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6990000000000000;

    #10 $display("\n1 * 2**665:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6980000000000000;

    #10 $display("\n1 * 2**664:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6970000000000000;

    #10 $display("\n1 * 2**663:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6960000000000000;

    #10 $display("\n1 * 2**662:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6950000000000000;

    #10 $display("\n1 * 2**661:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6940000000000000;

    #10 $display("\n1 * 2**660:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6930000000000000;

    #10 $display("\n1 * 2**659:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6920000000000000;

    #10 $display("\n1 * 2**658:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6910000000000000;

    #10 $display("\n1 * 2**657:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6900000000000000;

    #10 $display("\n1 * 2**656:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h68F0000000000000;

    #10 $display("\n1 * 2**655:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h68E0000000000000;

    #10 $display("\n1 * 2**654:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h68D0000000000000;

    #10 $display("\n1 * 2**653:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h68C0000000000000;

    #10 $display("\n1 * 2**652:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h68B0000000000000;

    #10 $display("\n1 * 2**651:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h68A0000000000000;

    #10 $display("\n1 * 2**650:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6890000000000000;

    #10 $display("\n1 * 2**649:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6880000000000000;

    #10 $display("\n1 * 2**648:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6870000000000000;

    #10 $display("\n1 * 2**647:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6860000000000000;

    #10 $display("\n1 * 2**646:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6850000000000000;

    #10 $display("\n1 * 2**645:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6840000000000000;

    #10 $display("\n1 * 2**644:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6830000000000000;

    #10 $display("\n1 * 2**643:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6820000000000000;

    #10 $display("\n1 * 2**642:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6810000000000000;

    #10 $display("\n1 * 2**641:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6800000000000000;

    #10 $display("\n1 * 2**640:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h67F0000000000000;

    #10 $display("\n1 * 2**639:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h67E0000000000000;

    #10 $display("\n1 * 2**638:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h67D0000000000000;

    #10 $display("\n1 * 2**637:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h67C0000000000000;

    #10 $display("\n1 * 2**636:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h67B0000000000000;

    #10 $display("\n1 * 2**635:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h67A0000000000000;

    #10 $display("\n1 * 2**634:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6790000000000000;

    #10 $display("\n1 * 2**633:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6780000000000000;

    #10 $display("\n1 * 2**632:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6770000000000000;

    #10 $display("\n1 * 2**631:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6760000000000000;

    #10 $display("\n1 * 2**630:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6750000000000000;

    #10 $display("\n1 * 2**629:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6740000000000000;

    #10 $display("\n1 * 2**628:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6730000000000000;

    #10 $display("\n1 * 2**627:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6720000000000000;

    #10 $display("\n1 * 2**626:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6710000000000000;

    #10 $display("\n1 * 2**625:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6700000000000000;

    #10 $display("\n1 * 2**624:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h66F0000000000000;

    #10 $display("\n1 * 2**623:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h66E0000000000000;

    #10 $display("\n1 * 2**622:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h66D0000000000000;

    #10 $display("\n1 * 2**621:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h66C0000000000000;

    #10 $display("\n1 * 2**620:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h66B0000000000000;

    #10 $display("\n1 * 2**619:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h66A0000000000000;

    #10 $display("\n1 * 2**618:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6690000000000000;

    #10 $display("\n1 * 2**617:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6680000000000000;

    #10 $display("\n1 * 2**616:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6670000000000000;

    #10 $display("\n1 * 2**615:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6660000000000000;

    #10 $display("\n1 * 2**614:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6650000000000000;

    #10 $display("\n1 * 2**613:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6640000000000000;

    #10 $display("\n1 * 2**612:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6630000000000000;

    #10 $display("\n1 * 2**611:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6620000000000000;

    #10 $display("\n1 * 2**610:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6610000000000000;

    #10 $display("\n1 * 2**609:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6600000000000000;

    #10 $display("\n1 * 2**608:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h65F0000000000000;

    #10 $display("\n1 * 2**607:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h65E0000000000000;

    #10 $display("\n1 * 2**606:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h65D0000000000000;

    #10 $display("\n1 * 2**605:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h65C0000000000000;

    #10 $display("\n1 * 2**604:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h65B0000000000000;

    #10 $display("\n1 * 2**603:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h65A0000000000000;

    #10 $display("\n1 * 2**602:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6590000000000000;

    #10 $display("\n1 * 2**601:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6580000000000000;

    #10 $display("\n1 * 2**600:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6570000000000000;

    #10 $display("\n1 * 2**599:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6560000000000000;

    #10 $display("\n1 * 2**598:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6550000000000000;

    #10 $display("\n1 * 2**597:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6540000000000000;

    #10 $display("\n1 * 2**596:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6530000000000000;

    #10 $display("\n1 * 2**595:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6520000000000000;

    #10 $display("\n1 * 2**594:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6510000000000000;

    #10 $display("\n1 * 2**593:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6500000000000000;

    #10 $display("\n1 * 2**592:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h64F0000000000000;

    #10 $display("\n1 * 2**591:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h64E0000000000000;

    #10 $display("\n1 * 2**590:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h64D0000000000000;

    #10 $display("\n1 * 2**589:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h64C0000000000000;

    #10 $display("\n1 * 2**588:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h64B0000000000000;

    #10 $display("\n1 * 2**587:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h64A0000000000000;

    #10 $display("\n1 * 2**586:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6490000000000000;

    #10 $display("\n1 * 2**585:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6480000000000000;

    #10 $display("\n1 * 2**584:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6470000000000000;

    #10 $display("\n1 * 2**583:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6460000000000000;

    #10 $display("\n1 * 2**582:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6450000000000000;

    #10 $display("\n1 * 2**581:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6440000000000000;

    #10 $display("\n1 * 2**580:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6430000000000000;

    #10 $display("\n1 * 2**579:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6420000000000000;

    #10 $display("\n1 * 2**578:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6410000000000000;

    #10 $display("\n1 * 2**577:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6400000000000000;

    #10 $display("\n1 * 2**576:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h63F0000000000000;

    #10 $display("\n1 * 2**575:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h63E0000000000000;

    #10 $display("\n1 * 2**574:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h63D0000000000000;

    #10 $display("\n1 * 2**573:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h63C0000000000000;

    #10 $display("\n1 * 2**572:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h63B0000000000000;

    #10 $display("\n1 * 2**571:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h63A0000000000000;

    #10 $display("\n1 * 2**570:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6390000000000000;

    #10 $display("\n1 * 2**569:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6380000000000000;

    #10 $display("\n1 * 2**568:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6370000000000000;

    #10 $display("\n1 * 2**567:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6360000000000000;

    #10 $display("\n1 * 2**566:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6350000000000000;

    #10 $display("\n1 * 2**565:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6340000000000000;

    #10 $display("\n1 * 2**564:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6330000000000000;

    #10 $display("\n1 * 2**563:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6320000000000000;

    #10 $display("\n1 * 2**562:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6310000000000000;

    #10 $display("\n1 * 2**561:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6300000000000000;

    #10 $display("\n1 * 2**560:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h62F0000000000000;

    #10 $display("\n1 * 2**559:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h62E0000000000000;

    #10 $display("\n1 * 2**558:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h62D0000000000000;

    #10 $display("\n1 * 2**557:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h62C0000000000000;

    #10 $display("\n1 * 2**556:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h62B0000000000000;

    #10 $display("\n1 * 2**555:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h62A0000000000000;

    #10 $display("\n1 * 2**554:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6290000000000000;

    #10 $display("\n1 * 2**553:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6280000000000000;

    #10 $display("\n1 * 2**552:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6270000000000000;

    #10 $display("\n1 * 2**551:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6260000000000000;

    #10 $display("\n1 * 2**550:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6250000000000000;

    #10 $display("\n1 * 2**549:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6240000000000000;

    #10 $display("\n1 * 2**548:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6230000000000000;

    #10 $display("\n1 * 2**547:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6220000000000000;

    #10 $display("\n1 * 2**546:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6210000000000000;

    #10 $display("\n1 * 2**545:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6200000000000000;

    #10 $display("\n1 * 2**544:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h61F0000000000000;

    #10 $display("\n1 * 2**543:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h61E0000000000000;

    #10 $display("\n1 * 2**542:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h61D0000000000000;

    #10 $display("\n1 * 2**541:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h61C0000000000000;

    #10 $display("\n1 * 2**540:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h61B0000000000000;

    #10 $display("\n1 * 2**539:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h61A0000000000000;

    #10 $display("\n1 * 2**538:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6190000000000000;

    #10 $display("\n1 * 2**537:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6180000000000000;

    #10 $display("\n1 * 2**536:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6170000000000000;

    #10 $display("\n1 * 2**535:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6160000000000000;

    #10 $display("\n1 * 2**534:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6150000000000000;

    #10 $display("\n1 * 2**533:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6140000000000000;

    #10 $display("\n1 * 2**532:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6130000000000000;

    #10 $display("\n1 * 2**531:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6120000000000000;

    #10 $display("\n1 * 2**530:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6110000000000000;

    #10 $display("\n1 * 2**529:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6100000000000000;

    #10 $display("\n1 * 2**528:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h60F0000000000000;

    #10 $display("\n1 * 2**527:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h60E0000000000000;

    #10 $display("\n1 * 2**526:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h60D0000000000000;

    #10 $display("\n1 * 2**525:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h60C0000000000000;

    #10 $display("\n1 * 2**524:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h60B0000000000000;

    #10 $display("\n1 * 2**523:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h60A0000000000000;

    #10 $display("\n1 * 2**522:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6090000000000000;

    #10 $display("\n1 * 2**521:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6080000000000000;

    #10 $display("\n1 * 2**520:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6070000000000000;

    #10 $display("\n1 * 2**519:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6060000000000000;

    #10 $display("\n1 * 2**518:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6050000000000000;

    #10 $display("\n1 * 2**517:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6040000000000000;

    #10 $display("\n1 * 2**516:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6030000000000000;

    #10 $display("\n1 * 2**515:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6020000000000000;

    #10 $display("\n1 * 2**514:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6010000000000000;

    #10 $display("\n1 * 2**513:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h6000000000000000;

    #10 $display("\n1 * 2**512:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5FF0000000000000;

    #10 $display("\n1 * 2**511:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5FE0000000000000;

    #10 $display("\n1 * 2**510:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5FD0000000000000;

    #10 $display("\n1 * 2**509:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5FC0000000000000;

    #10 $display("\n1 * 2**508:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5FB0000000000000;

    #10 $display("\n1 * 2**507:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5FA0000000000000;

    #10 $display("\n1 * 2**506:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5F90000000000000;

    #10 $display("\n1 * 2**505:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5F80000000000000;

    #10 $display("\n1 * 2**504:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5F70000000000000;

    #10 $display("\n1 * 2**503:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5F60000000000000;

    #10 $display("\n1 * 2**502:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5F50000000000000;

    #10 $display("\n1 * 2**501:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5F40000000000000;

    #10 $display("\n1 * 2**500:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5F30000000000000;

    #10 $display("\n1 * 2**499:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5F20000000000000;

    #10 $display("\n1 * 2**498:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5F10000000000000;

    #10 $display("\n1 * 2**497:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5F00000000000000;

    #10 $display("\n1 * 2**496:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5EF0000000000000;

    #10 $display("\n1 * 2**495:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5EE0000000000000;

    #10 $display("\n1 * 2**494:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5ED0000000000000;

    #10 $display("\n1 * 2**493:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5EC0000000000000;

    #10 $display("\n1 * 2**492:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5EB0000000000000;

    #10 $display("\n1 * 2**491:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5EA0000000000000;

    #10 $display("\n1 * 2**490:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5E90000000000000;

    #10 $display("\n1 * 2**489:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5E80000000000000;

    #10 $display("\n1 * 2**488:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5E70000000000000;

    #10 $display("\n1 * 2**487:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5E60000000000000;

    #10 $display("\n1 * 2**486:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5E50000000000000;

    #10 $display("\n1 * 2**485:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5E40000000000000;

    #10 $display("\n1 * 2**484:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5E30000000000000;

    #10 $display("\n1 * 2**483:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5E20000000000000;

    #10 $display("\n1 * 2**482:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5E10000000000000;

    #10 $display("\n1 * 2**481:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5E00000000000000;

    #10 $display("\n1 * 2**480:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5DF0000000000000;

    #10 $display("\n1 * 2**479:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5DE0000000000000;

    #10 $display("\n1 * 2**478:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5DD0000000000000;

    #10 $display("\n1 * 2**477:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5DC0000000000000;

    #10 $display("\n1 * 2**476:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5DB0000000000000;

    #10 $display("\n1 * 2**475:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5DA0000000000000;

    #10 $display("\n1 * 2**474:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5D90000000000000;

    #10 $display("\n1 * 2**473:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5D80000000000000;

    #10 $display("\n1 * 2**472:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5D70000000000000;

    #10 $display("\n1 * 2**471:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5D60000000000000;

    #10 $display("\n1 * 2**470:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5D50000000000000;

    #10 $display("\n1 * 2**469:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5D40000000000000;

    #10 $display("\n1 * 2**468:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5D30000000000000;

    #10 $display("\n1 * 2**467:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5D20000000000000;

    #10 $display("\n1 * 2**466:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5D10000000000000;

    #10 $display("\n1 * 2**465:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5D00000000000000;

    #10 $display("\n1 * 2**464:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5CF0000000000000;

    #10 $display("\n1 * 2**463:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5CE0000000000000;

    #10 $display("\n1 * 2**462:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5CD0000000000000;

    #10 $display("\n1 * 2**461:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5CC0000000000000;

    #10 $display("\n1 * 2**460:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5CB0000000000000;

    #10 $display("\n1 * 2**459:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5CA0000000000000;

    #10 $display("\n1 * 2**458:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5C90000000000000;

    #10 $display("\n1 * 2**457:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5C80000000000000;

    #10 $display("\n1 * 2**456:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5C70000000000000;

    #10 $display("\n1 * 2**455:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5C60000000000000;

    #10 $display("\n1 * 2**454:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5C50000000000000;

    #10 $display("\n1 * 2**453:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5C40000000000000;

    #10 $display("\n1 * 2**452:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5C30000000000000;

    #10 $display("\n1 * 2**451:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5C20000000000000;

    #10 $display("\n1 * 2**450:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5C10000000000000;

    #10 $display("\n1 * 2**449:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5C00000000000000;

    #10 $display("\n1 * 2**448:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5BF0000000000000;

    #10 $display("\n1 * 2**447:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5BE0000000000000;

    #10 $display("\n1 * 2**446:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5BD0000000000000;

    #10 $display("\n1 * 2**445:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5BC0000000000000;

    #10 $display("\n1 * 2**444:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5BB0000000000000;

    #10 $display("\n1 * 2**443:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5BA0000000000000;

    #10 $display("\n1 * 2**442:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5B90000000000000;

    #10 $display("\n1 * 2**441:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5B80000000000000;

    #10 $display("\n1 * 2**440:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5B70000000000000;

    #10 $display("\n1 * 2**439:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5B60000000000000;

    #10 $display("\n1 * 2**438:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5B50000000000000;

    #10 $display("\n1 * 2**437:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5B40000000000000;

    #10 $display("\n1 * 2**436:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5B30000000000000;

    #10 $display("\n1 * 2**435:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5B20000000000000;

    #10 $display("\n1 * 2**434:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5B10000000000000;

    #10 $display("\n1 * 2**433:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5B00000000000000;

    #10 $display("\n1 * 2**432:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5AF0000000000000;

    #10 $display("\n1 * 2**431:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5AE0000000000000;

    #10 $display("\n1 * 2**430:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5AD0000000000000;

    #10 $display("\n1 * 2**429:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5AC0000000000000;

    #10 $display("\n1 * 2**428:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5AB0000000000000;

    #10 $display("\n1 * 2**427:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5AA0000000000000;

    #10 $display("\n1 * 2**426:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5A90000000000000;

    #10 $display("\n1 * 2**425:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5A80000000000000;

    #10 $display("\n1 * 2**424:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5A70000000000000;

    #10 $display("\n1 * 2**423:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5A60000000000000;

    #10 $display("\n1 * 2**422:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5A50000000000000;

    #10 $display("\n1 * 2**421:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5A40000000000000;

    #10 $display("\n1 * 2**420:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5A30000000000000;

    #10 $display("\n1 * 2**419:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5A20000000000000;

    #10 $display("\n1 * 2**418:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5A10000000000000;

    #10 $display("\n1 * 2**417:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5A00000000000000;

    #10 $display("\n1 * 2**416:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h59F0000000000000;

    #10 $display("\n1 * 2**415:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h59E0000000000000;

    #10 $display("\n1 * 2**414:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h59D0000000000000;

    #10 $display("\n1 * 2**413:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h59C0000000000000;

    #10 $display("\n1 * 2**412:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h59B0000000000000;

    #10 $display("\n1 * 2**411:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h59A0000000000000;

    #10 $display("\n1 * 2**410:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5990000000000000;

    #10 $display("\n1 * 2**409:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5980000000000000;

    #10 $display("\n1 * 2**408:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5970000000000000;

    #10 $display("\n1 * 2**407:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5960000000000000;

    #10 $display("\n1 * 2**406:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5950000000000000;

    #10 $display("\n1 * 2**405:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5940000000000000;

    #10 $display("\n1 * 2**404:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5930000000000000;

    #10 $display("\n1 * 2**403:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5920000000000000;

    #10 $display("\n1 * 2**402:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5910000000000000;

    #10 $display("\n1 * 2**401:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5900000000000000;

    #10 $display("\n1 * 2**400:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h58F0000000000000;

    #10 $display("\n1 * 2**399:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h58E0000000000000;

    #10 $display("\n1 * 2**398:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h58D0000000000000;

    #10 $display("\n1 * 2**397:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h58C0000000000000;

    #10 $display("\n1 * 2**396:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h58B0000000000000;

    #10 $display("\n1 * 2**395:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h58A0000000000000;

    #10 $display("\n1 * 2**394:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5890000000000000;

    #10 $display("\n1 * 2**393:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5880000000000000;

    #10 $display("\n1 * 2**392:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5870000000000000;

    #10 $display("\n1 * 2**391:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5860000000000000;

    #10 $display("\n1 * 2**390:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5850000000000000;

    #10 $display("\n1 * 2**389:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5840000000000000;

    #10 $display("\n1 * 2**388:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5830000000000000;

    #10 $display("\n1 * 2**387:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5820000000000000;

    #10 $display("\n1 * 2**386:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5810000000000000;

    #10 $display("\n1 * 2**385:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5800000000000000;

    #10 $display("\n1 * 2**384:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h57F0000000000000;

    #10 $display("\n1 * 2**383:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h57E0000000000000;

    #10 $display("\n1 * 2**382:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h57D0000000000000;

    #10 $display("\n1 * 2**381:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h57C0000000000000;

    #10 $display("\n1 * 2**380:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h57B0000000000000;

    #10 $display("\n1 * 2**379:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h57A0000000000000;

    #10 $display("\n1 * 2**378:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5790000000000000;

    #10 $display("\n1 * 2**377:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5780000000000000;

    #10 $display("\n1 * 2**376:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5770000000000000;

    #10 $display("\n1 * 2**375:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5760000000000000;

    #10 $display("\n1 * 2**374:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5750000000000000;

    #10 $display("\n1 * 2**373:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5740000000000000;

    #10 $display("\n1 * 2**372:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5730000000000000;

    #10 $display("\n1 * 2**371:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5720000000000000;

    #10 $display("\n1 * 2**370:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5710000000000000;

    #10 $display("\n1 * 2**369:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5700000000000000;

    #10 $display("\n1 * 2**368:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h56F0000000000000;

    #10 $display("\n1 * 2**367:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h56E0000000000000;

    #10 $display("\n1 * 2**366:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h56D0000000000000;

    #10 $display("\n1 * 2**365:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h56C0000000000000;

    #10 $display("\n1 * 2**364:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h56B0000000000000;

    #10 $display("\n1 * 2**363:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h56A0000000000000;

    #10 $display("\n1 * 2**362:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5690000000000000;

    #10 $display("\n1 * 2**361:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5680000000000000;

    #10 $display("\n1 * 2**360:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5670000000000000;

    #10 $display("\n1 * 2**359:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5660000000000000;

    #10 $display("\n1 * 2**358:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5650000000000000;

    #10 $display("\n1 * 2**357:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5640000000000000;

    #10 $display("\n1 * 2**356:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5630000000000000;

    #10 $display("\n1 * 2**355:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5620000000000000;

    #10 $display("\n1 * 2**354:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5610000000000000;

    #10 $display("\n1 * 2**353:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5600000000000000;

    #10 $display("\n1 * 2**352:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h55F0000000000000;

    #10 $display("\n1 * 2**351:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h55E0000000000000;

    #10 $display("\n1 * 2**350:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h55D0000000000000;

    #10 $display("\n1 * 2**349:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h55C0000000000000;

    #10 $display("\n1 * 2**348:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h55B0000000000000;

    #10 $display("\n1 * 2**347:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h55A0000000000000;

    #10 $display("\n1 * 2**346:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5590000000000000;

    #10 $display("\n1 * 2**345:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5580000000000000;

    #10 $display("\n1 * 2**344:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5570000000000000;

    #10 $display("\n1 * 2**343:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5560000000000000;

    #10 $display("\n1 * 2**342:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5550000000000000;

    #10 $display("\n1 * 2**341:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5540000000000000;

    #10 $display("\n1 * 2**340:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5530000000000000;

    #10 $display("\n1 * 2**339:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5520000000000000;

    #10 $display("\n1 * 2**338:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5510000000000000;

    #10 $display("\n1 * 2**337:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5500000000000000;

    #10 $display("\n1 * 2**336:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h54F0000000000000;

    #10 $display("\n1 * 2**335:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h54E0000000000000;

    #10 $display("\n1 * 2**334:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h54D0000000000000;

    #10 $display("\n1 * 2**333:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h54C0000000000000;

    #10 $display("\n1 * 2**332:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h54B0000000000000;

    #10 $display("\n1 * 2**331:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h54A0000000000000;

    #10 $display("\n1 * 2**330:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5490000000000000;

    #10 $display("\n1 * 2**329:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5480000000000000;

    #10 $display("\n1 * 2**328:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5470000000000000;

    #10 $display("\n1 * 2**327:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5460000000000000;

    #10 $display("\n1 * 2**326:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5450000000000000;

    #10 $display("\n1 * 2**325:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5440000000000000;

    #10 $display("\n1 * 2**324:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5430000000000000;

    #10 $display("\n1 * 2**323:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5420000000000000;

    #10 $display("\n1 * 2**322:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5410000000000000;

    #10 $display("\n1 * 2**321:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5400000000000000;

    #10 $display("\n1 * 2**320:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h53F0000000000000;

    #10 $display("\n1 * 2**319:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h53E0000000000000;

    #10 $display("\n1 * 2**318:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h53D0000000000000;

    #10 $display("\n1 * 2**317:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h53C0000000000000;

    #10 $display("\n1 * 2**316:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h53B0000000000000;

    #10 $display("\n1 * 2**315:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h53A0000000000000;

    #10 $display("\n1 * 2**314:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5390000000000000;

    #10 $display("\n1 * 2**313:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5380000000000000;

    #10 $display("\n1 * 2**312:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5370000000000000;

    #10 $display("\n1 * 2**311:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5360000000000000;

    #10 $display("\n1 * 2**310:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5350000000000000;

    #10 $display("\n1 * 2**309:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5340000000000000;

    #10 $display("\n1 * 2**308:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5330000000000000;

    #10 $display("\n1 * 2**307:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5320000000000000;

    #10 $display("\n1 * 2**306:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5310000000000000;

    #10 $display("\n1 * 2**305:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5300000000000000;

    #10 $display("\n1 * 2**304:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h52F0000000000000;

    #10 $display("\n1 * 2**303:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h52E0000000000000;

    #10 $display("\n1 * 2**302:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h52D0000000000000;

    #10 $display("\n1 * 2**301:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h52C0000000000000;

    #10 $display("\n1 * 2**300:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h52B0000000000000;

    #10 $display("\n1 * 2**299:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h52A0000000000000;

    #10 $display("\n1 * 2**298:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5290000000000000;

    #10 $display("\n1 * 2**297:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5280000000000000;

    #10 $display("\n1 * 2**296:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5270000000000000;

    #10 $display("\n1 * 2**295:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5260000000000000;

    #10 $display("\n1 * 2**294:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5250000000000000;

    #10 $display("\n1 * 2**293:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5240000000000000;

    #10 $display("\n1 * 2**292:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5230000000000000;

    #10 $display("\n1 * 2**291:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5220000000000000;

    #10 $display("\n1 * 2**290:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5210000000000000;

    #10 $display("\n1 * 2**289:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5200000000000000;

    #10 $display("\n1 * 2**288:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h51F0000000000000;

    #10 $display("\n1 * 2**287:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h51E0000000000000;

    #10 $display("\n1 * 2**286:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h51D0000000000000;

    #10 $display("\n1 * 2**285:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h51C0000000000000;

    #10 $display("\n1 * 2**284:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h51B0000000000000;

    #10 $display("\n1 * 2**283:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h51A0000000000000;

    #10 $display("\n1 * 2**282:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5190000000000000;

    #10 $display("\n1 * 2**281:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5180000000000000;

    #10 $display("\n1 * 2**280:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5170000000000000;

    #10 $display("\n1 * 2**279:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5160000000000000;

    #10 $display("\n1 * 2**278:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5150000000000000;

    #10 $display("\n1 * 2**277:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5140000000000000;

    #10 $display("\n1 * 2**276:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5130000000000000;

    #10 $display("\n1 * 2**275:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5120000000000000;

    #10 $display("\n1 * 2**274:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5110000000000000;

    #10 $display("\n1 * 2**273:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5100000000000000;

    #10 $display("\n1 * 2**272:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h50F0000000000000;

    #10 $display("\n1 * 2**271:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h50E0000000000000;

    #10 $display("\n1 * 2**270:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h50D0000000000000;

    #10 $display("\n1 * 2**269:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h50C0000000000000;

    #10 $display("\n1 * 2**268:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h50B0000000000000;

    #10 $display("\n1 * 2**267:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h50A0000000000000;

    #10 $display("\n1 * 2**266:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5090000000000000;

    #10 $display("\n1 * 2**265:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5080000000000000;

    #10 $display("\n1 * 2**264:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5070000000000000;

    #10 $display("\n1 * 2**263:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5060000000000000;

    #10 $display("\n1 * 2**262:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5050000000000000;

    #10 $display("\n1 * 2**261:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5040000000000000;

    #10 $display("\n1 * 2**260:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5030000000000000;

    #10 $display("\n1 * 2**259:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5020000000000000;

    #10 $display("\n1 * 2**258:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5010000000000000;

    #10 $display("\n1 * 2**257:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h5000000000000000;

    #10 $display("\n1 * 2**256:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4FF0000000000000;

    #10 $display("\n1 * 2**255:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4FE0000000000000;

    #10 $display("\n1 * 2**254:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4FD0000000000000;

    #10 $display("\n1 * 2**253:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4FC0000000000000;

    #10 $display("\n1 * 2**252:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4FB0000000000000;

    #10 $display("\n1 * 2**251:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4FA0000000000000;

    #10 $display("\n1 * 2**250:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4F90000000000000;

    #10 $display("\n1 * 2**249:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4F80000000000000;

    #10 $display("\n1 * 2**248:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4F70000000000000;

    #10 $display("\n1 * 2**247:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4F60000000000000;

    #10 $display("\n1 * 2**246:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4F50000000000000;

    #10 $display("\n1 * 2**245:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4F40000000000000;

    #10 $display("\n1 * 2**244:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4F30000000000000;

    #10 $display("\n1 * 2**243:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4F20000000000000;

    #10 $display("\n1 * 2**242:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4F10000000000000;

    #10 $display("\n1 * 2**241:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4F00000000000000;

    #10 $display("\n1 * 2**240:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4EF0000000000000;

    #10 $display("\n1 * 2**239:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4EE0000000000000;

    #10 $display("\n1 * 2**238:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4ED0000000000000;

    #10 $display("\n1 * 2**237:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4EC0000000000000;

    #10 $display("\n1 * 2**236:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4EB0000000000000;

    #10 $display("\n1 * 2**235:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4EA0000000000000;

    #10 $display("\n1 * 2**234:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4E90000000000000;

    #10 $display("\n1 * 2**233:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4E80000000000000;

    #10 $display("\n1 * 2**232:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4E70000000000000;

    #10 $display("\n1 * 2**231:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4E60000000000000;

    #10 $display("\n1 * 2**230:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4E50000000000000;

    #10 $display("\n1 * 2**229:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4E40000000000000;

    #10 $display("\n1 * 2**228:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4E30000000000000;

    #10 $display("\n1 * 2**227:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4E20000000000000;

    #10 $display("\n1 * 2**226:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4E10000000000000;

    #10 $display("\n1 * 2**225:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4E00000000000000;

    #10 $display("\n1 * 2**224:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4DF0000000000000;

    #10 $display("\n1 * 2**223:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4DE0000000000000;

    #10 $display("\n1 * 2**222:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4DD0000000000000;

    #10 $display("\n1 * 2**221:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4DC0000000000000;

    #10 $display("\n1 * 2**220:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4DB0000000000000;

    #10 $display("\n1 * 2**219:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4DA0000000000000;

    #10 $display("\n1 * 2**218:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4D90000000000000;

    #10 $display("\n1 * 2**217:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4D80000000000000;

    #10 $display("\n1 * 2**216:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4D70000000000000;

    #10 $display("\n1 * 2**215:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4D60000000000000;

    #10 $display("\n1 * 2**214:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4D50000000000000;

    #10 $display("\n1 * 2**213:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4D40000000000000;

    #10 $display("\n1 * 2**212:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4D30000000000000;

    #10 $display("\n1 * 2**211:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4D20000000000000;

    #10 $display("\n1 * 2**210:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4D10000000000000;

    #10 $display("\n1 * 2**209:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4D00000000000000;

    #10 $display("\n1 * 2**208:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4CF0000000000000;

    #10 $display("\n1 * 2**207:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4CE0000000000000;

    #10 $display("\n1 * 2**206:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4CD0000000000000;

    #10 $display("\n1 * 2**205:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4CC0000000000000;

    #10 $display("\n1 * 2**204:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4CB0000000000000;

    #10 $display("\n1 * 2**203:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4CA0000000000000;

    #10 $display("\n1 * 2**202:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4C90000000000000;

    #10 $display("\n1 * 2**201:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4C80000000000000;

    #10 $display("\n1 * 2**200:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4C70000000000000;

    #10 $display("\n1 * 2**199:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4C60000000000000;

    #10 $display("\n1 * 2**198:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4C50000000000000;

    #10 $display("\n1 * 2**197:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4C40000000000000;

    #10 $display("\n1 * 2**196:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4C30000000000000;

    #10 $display("\n1 * 2**195:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4C20000000000000;

    #10 $display("\n1 * 2**194:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4C10000000000000;

    #10 $display("\n1 * 2**193:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4C00000000000000;

    #10 $display("\n1 * 2**192:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4BF0000000000000;

    #10 $display("\n1 * 2**191:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4BE0000000000000;

    #10 $display("\n1 * 2**190:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4BD0000000000000;

    #10 $display("\n1 * 2**189:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4BC0000000000000;

    #10 $display("\n1 * 2**188:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4BB0000000000000;

    #10 $display("\n1 * 2**187:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4BA0000000000000;

    #10 $display("\n1 * 2**186:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4B90000000000000;

    #10 $display("\n1 * 2**185:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4B80000000000000;

    #10 $display("\n1 * 2**184:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4B70000000000000;

    #10 $display("\n1 * 2**183:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4B60000000000000;

    #10 $display("\n1 * 2**182:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4B50000000000000;

    #10 $display("\n1 * 2**181:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4B40000000000000;

    #10 $display("\n1 * 2**180:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4B30000000000000;

    #10 $display("\n1 * 2**179:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4B20000000000000;

    #10 $display("\n1 * 2**178:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4B10000000000000;

    #10 $display("\n1 * 2**177:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4B00000000000000;

    #10 $display("\n1 * 2**176:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4AF0000000000000;

    #10 $display("\n1 * 2**175:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4AE0000000000000;

    #10 $display("\n1 * 2**174:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4AD0000000000000;

    #10 $display("\n1 * 2**173:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4AC0000000000000;

    #10 $display("\n1 * 2**172:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4AB0000000000000;

    #10 $display("\n1 * 2**171:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4AA0000000000000;

    #10 $display("\n1 * 2**170:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4A90000000000000;

    #10 $display("\n1 * 2**169:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4A80000000000000;

    #10 $display("\n1 * 2**168:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4A70000000000000;

    #10 $display("\n1 * 2**167:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4A60000000000000;

    #10 $display("\n1 * 2**166:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4A50000000000000;

    #10 $display("\n1 * 2**165:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4A40000000000000;

    #10 $display("\n1 * 2**164:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4A30000000000000;

    #10 $display("\n1 * 2**163:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4A20000000000000;

    #10 $display("\n1 * 2**162:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4A10000000000000;

    #10 $display("\n1 * 2**161:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4A00000000000000;

    #10 $display("\n1 * 2**160:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h49F0000000000000;

    #10 $display("\n1 * 2**159:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h49E0000000000000;

    #10 $display("\n1 * 2**158:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h49D0000000000000;

    #10 $display("\n1 * 2**157:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h49C0000000000000;

    #10 $display("\n1 * 2**156:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h49B0000000000000;

    #10 $display("\n1 * 2**155:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h49A0000000000000;

    #10 $display("\n1 * 2**154:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4990000000000000;

    #10 $display("\n1 * 2**153:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4980000000000000;

    #10 $display("\n1 * 2**152:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4970000000000000;

    #10 $display("\n1 * 2**151:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4960000000000000;

    #10 $display("\n1 * 2**150:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4950000000000000;

    #10 $display("\n1 * 2**149:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4940000000000000;

    #10 $display("\n1 * 2**148:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4930000000000000;

    #10 $display("\n1 * 2**147:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4920000000000000;

    #10 $display("\n1 * 2**146:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4910000000000000;

    #10 $display("\n1 * 2**145:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4900000000000000;

    #10 $display("\n1 * 2**144:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h48F0000000000000;

    #10 $display("\n1 * 2**143:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h48E0000000000000;

    #10 $display("\n1 * 2**142:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h48D0000000000000;

    #10 $display("\n1 * 2**141:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h48C0000000000000;

    #10 $display("\n1 * 2**140:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h48B0000000000000;

    #10 $display("\n1 * 2**139:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h48A0000000000000;

    #10 $display("\n1 * 2**138:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4890000000000000;

    #10 $display("\n1 * 2**137:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4880000000000000;

    #10 $display("\n1 * 2**136:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4870000000000000;

    #10 $display("\n1 * 2**135:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4860000000000000;

    #10 $display("\n1 * 2**134:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4850000000000000;

    #10 $display("\n1 * 2**133:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4840000000000000;

    #10 $display("\n1 * 2**132:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4830000000000000;

    #10 $display("\n1 * 2**131:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4820000000000000;

    #10 $display("\n1 * 2**130:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4810000000000000;

    #10 $display("\n1 * 2**129:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4800000000000000;

    #10 $display("\n1 * 2**128:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h47F0000000000000;

    #10 $display("\n1 * 2**127:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h47E0000000000000;

    #10 $display("\n1 * 2**126:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h47D0000000000000;

    #10 $display("\n1 * 2**125:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h47C0000000000000;

    #10 $display("\n1 * 2**124:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h47B0000000000000;

    #10 $display("\n1 * 2**123:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h47A0000000000000;

    #10 $display("\n1 * 2**122:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4790000000000000;

    #10 $display("\n1 * 2**121:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4780000000000000;

    #10 $display("\n1 * 2**120:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4770000000000000;

    #10 $display("\n1 * 2**119:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4760000000000000;

    #10 $display("\n1 * 2**118:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4750000000000000;

    #10 $display("\n1 * 2**117:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4740000000000000;

    #10 $display("\n1 * 2**116:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4730000000000000;

    #10 $display("\n1 * 2**115:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4720000000000000;

    #10 $display("\n1 * 2**114:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4710000000000000;

    #10 $display("\n1 * 2**113:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4700000000000000;

    #10 $display("\n1 * 2**112:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h46F0000000000000;

    #10 $display("\n1 * 2**111:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h46E0000000000000;

    #10 $display("\n1 * 2**110:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h46D0000000000000;

    #10 $display("\n1 * 2**109:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h46C0000000000000;

    #10 $display("\n1 * 2**108:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h46B0000000000000;

    #10 $display("\n1 * 2**107:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h46A0000000000000;

    #10 $display("\n1 * 2**106:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4690000000000000;

    #10 $display("\n1 * 2**105:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4680000000000000;

    #10 $display("\n1 * 2**104:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4670000000000000;

    #10 $display("\n1 * 2**103:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4660000000000000;

    #10 $display("\n1 * 2**102:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4650000000000000;

    #10 $display("\n1 * 2**101:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4640000000000000;

    #10 $display("\n1 * 2**100:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4630000000000000;

    #10 $display("\n1 * 2**99:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4620000000000000;

    #10 $display("\n1 * 2**98:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4610000000000000;

    #10 $display("\n1 * 2**97:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4600000000000000;

    #10 $display("\n1 * 2**96:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h45F0000000000000;

    #10 $display("\n1 * 2**95:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h45E0000000000000;

    #10 $display("\n1 * 2**94:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h45D0000000000000;

    #10 $display("\n1 * 2**93:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h45C0000000000000;

    #10 $display("\n1 * 2**92:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h45B0000000000000;

    #10 $display("\n1 * 2**91:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h45A0000000000000;

    #10 $display("\n1 * 2**90:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4590000000000000;

    #10 $display("\n1 * 2**89:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4580000000000000;

    #10 $display("\n1 * 2**88:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4570000000000000;

    #10 $display("\n1 * 2**87:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4560000000000000;

    #10 $display("\n1 * 2**86:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4550000000000000;

    #10 $display("\n1 * 2**85:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4540000000000000;

    #10 $display("\n1 * 2**84:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4530000000000000;

    #10 $display("\n1 * 2**83:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4520000000000000;

    #10 $display("\n1 * 2**82:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4510000000000000;

    #10 $display("\n1 * 2**81:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4500000000000000;

    #10 $display("\n1 * 2**80:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h44F0000000000000;

    #10 $display("\n1 * 2**79:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h44E0000000000000;

    #10 $display("\n1 * 2**78:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h44D0000000000000;

    #10 $display("\n1 * 2**77:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h44C0000000000000;

    #10 $display("\n1 * 2**76:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h44B0000000000000;

    #10 $display("\n1 * 2**75:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h44A0000000000000;

    #10 $display("\n1 * 2**74:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4490000000000000;

    #10 $display("\n1 * 2**73:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4480000000000000;

    #10 $display("\n1 * 2**72:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4470000000000000;

    #10 $display("\n1 * 2**71:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4460000000000000;

    #10 $display("\n1 * 2**70:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4450000000000000;

    #10 $display("\n1 * 2**69:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4440000000000000;

    #10 $display("\n1 * 2**68:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4430000000000000;

    #10 $display("\n1 * 2**67:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4420000000000000;

    #10 $display("\n1 * 2**66:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4410000000000000;

    #10 $display("\n1 * 2**65:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4400000000000000;

    #10 $display("\n1 * 2**64:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h43F0000000000000;

    #10 $display("\n1 * 2**63:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h43E0000000000000;

    #10 $display("\n1 * 2**62:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h43D0000000000000;

    #10 $display("\n1 * 2**61:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h43C0000000000000;

    #10 $display("\n1 * 2**60:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h43B0000000000000;

    #10 $display("\n1 * 2**59:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h43A0000000000000;

    #10 $display("\n1 * 2**58:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4390000000000000;

    #10 $display("\n1 * 2**57:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4380000000000000;

    #10 $display("\n1 * 2**56:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4370000000000000;

    #10 $display("\n1 * 2**55:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4360000000000000;

    #10 $display("\n1 * 2**54:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4350000000000000;

    #10 $display("\n1 * 2**53:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4340000000000000;

    #10 $display("\n1 * 2**52:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4330000000000000;

    #10 $display("\n1 * 2**51:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4320000000000000;

    #10 $display("\n1 * 2**50:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4310000000000000;

    #10 $display("\n1 * 2**49:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4300000000000000;

    #10 $display("\n1 * 2**48:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h42F0000000000000;

    #10 $display("\n1 * 2**47:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h42E0000000000000;

    #10 $display("\n1 * 2**46:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h42D0000000000000;

    #10 $display("\n1 * 2**45:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h42C0000000000000;

    #10 $display("\n1 * 2**44:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h42B0000000000000;

    #10 $display("\n1 * 2**43:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h42A0000000000000;

    #10 $display("\n1 * 2**42:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4290000000000000;

    #10 $display("\n1 * 2**41:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4280000000000000;

    #10 $display("\n1 * 2**40:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4270000000000000;

    #10 $display("\n1 * 2**39:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4260000000000000;

    #10 $display("\n1 * 2**38:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4250000000000000;

    #10 $display("\n1 * 2**37:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4240000000000000;

    #10 $display("\n1 * 2**36:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4230000000000000;

    #10 $display("\n1 * 2**35:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4220000000000000;

    #10 $display("\n1 * 2**34:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4210000000000000;

    #10 $display("\n1 * 2**33:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4200000000000000;

    #10 $display("\n1 * 2**32:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h41F0000000000000;

    #10 $display("\n1 * 2**31:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h41E0000000000000;

    #10 $display("\n1 * 2**30:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h41D0000000000000;

    #10 $display("\n1 * 2**29:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h41C0000000000000;

    #10 $display("\n1 * 2**28:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h41B0000000000000;

    #10 $display("\n1 * 2**27:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h41A0000000000000;

    #10 $display("\n1 * 2**26:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4190000000000000;

    #10 $display("\n1 * 2**25:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4180000000000000;

    #10 $display("\n1 * 2**24:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4170000000000000;

    #10 $display("\n1 * 2**23:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4160000000000000;

    #10 $display("\n1 * 2**22:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4150000000000000;

    #10 $display("\n1 * 2**21:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4140000000000000;

    #10 $display("\n1 * 2**20:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4130000000000000;

    #10 $display("\n1 * 2**19:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4120000000000000;

    #10 $display("\n1 * 2**18:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4110000000000000;

    #10 $display("\n1 * 2**17:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4100000000000000;

    #10 $display("\n1 * 2**16:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h40F0000000000000;

    #10 $display("\n1 * 2**15:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h40E0000000000000;

    #10 $display("\n1 * 2**14:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h40D0000000000000;

    #10 $display("\n1 * 2**13:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h40C0000000000000;

    #10 $display("\n1 * 2**12:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h40B0000000000000;

    #10 $display("\n1 * 2**11:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h40A0000000000000;

    #10 $display("\n1 * 2**10:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4090000000000000;

    #10 $display("\n1 * 2**9:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4080000000000000;

    #10 $display("\n1 * 2**8:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4070000000000000;

    #10 $display("\n1 * 2**7:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4060000000000000;

    #10 $display("\n1 * 2**6:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4050000000000000;

    #10 $display("\n1 * 2**5:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4040000000000000;

    #10 $display("\n1 * 2**4:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4030000000000000;

    #10 $display("\n1 * 2**3:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4020000000000000;

    #10 $display("\n1 * 2**2:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4010000000000000;

    #10 $display("\n1 * 2**1:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h4000000000000000;

    #10 $display("\n1 * 2**0:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3FF0000000000000;

    #10 $display("\n1 * 2**-1:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3FE0000000000000;

    #10 $display("\n1 * 2**-2:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3FD0000000000000;

    #10 $display("\n1 * 2**-3:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3FC0000000000000;

    #10 $display("\n1 * 2**-4:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3FB0000000000000;

    #10 $display("\n1 * 2**-5:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3FA0000000000000;

    #10 $display("\n1 * 2**-6:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3F90000000000000;

    #10 $display("\n1 * 2**-7:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3F80000000000000;

    #10 $display("\n1 * 2**-8:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3F70000000000000;

    #10 $display("\n1 * 2**-9:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3F60000000000000;

    #10 $display("\n1 * 2**-10:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3F50000000000000;

    #10 $display("\n1 * 2**-11:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3F40000000000000;

    #10 $display("\n1 * 2**-12:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3F30000000000000;

    #10 $display("\n1 * 2**-13:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3F20000000000000;

    #10 $display("\n1 * 2**-14:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3F10000000000000;

    #10 $display("\n1 * 2**-15:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3F00000000000000;

    #10 $display("\n1 * 2**-16:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3EF0000000000000;

    #10 $display("\n1 * 2**-17:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3EE0000000000000;

    #10 $display("\n1 * 2**-18:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3ED0000000000000;

    #10 $display("\n1 * 2**-19:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3EC0000000000000;

    #10 $display("\n1 * 2**-20:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3EB0000000000000;

    #10 $display("\n1 * 2**-21:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3EA0000000000000;

    #10 $display("\n1 * 2**-22:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3E90000000000000;

    #10 $display("\n1 * 2**-23:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3E80000000000000;

    #10 $display("\n1 * 2**-24:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3E70000000000000;

    #10 $display("\n1 * 2**-25:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3E60000000000000;

    #10 $display("\n1 * 2**-26:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3E50000000000000;

    #10 $display("\n1 * 2**-27:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3E40000000000000;

    #10 $display("\n1 * 2**-28:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3E30000000000000;

    #10 $display("\n1 * 2**-29:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3E20000000000000;

    #10 $display("\n1 * 2**-30:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3E10000000000000;

    #10 $display("\n1 * 2**-31:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3E00000000000000;

    #10 $display("\n1 * 2**-32:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3DF0000000000000;

    #10 $display("\n1 * 2**-33:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3DE0000000000000;

    #10 $display("\n1 * 2**-34:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3DD0000000000000;

    #10 $display("\n1 * 2**-35:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3DC0000000000000;

    #10 $display("\n1 * 2**-36:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3DB0000000000000;

    #10 $display("\n1 * 2**-37:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3DA0000000000000;

    #10 $display("\n1 * 2**-38:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3D90000000000000;

    #10 $display("\n1 * 2**-39:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3D80000000000000;

    #10 $display("\n1 * 2**-40:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3D70000000000000;

    #10 $display("\n1 * 2**-41:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3D60000000000000;

    #10 $display("\n1 * 2**-42:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3D50000000000000;

    #10 $display("\n1 * 2**-43:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3D40000000000000;

    #10 $display("\n1 * 2**-44:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3D30000000000000;

    #10 $display("\n1 * 2**-45:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3D20000000000000;

    #10 $display("\n1 * 2**-46:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3D10000000000000;

    #10 $display("\n1 * 2**-47:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3D00000000000000;

    #10 $display("\n1 * 2**-48:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3CF0000000000000;

    #10 $display("\n1 * 2**-49:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3CE0000000000000;

    #10 $display("\n1 * 2**-50:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3CD0000000000000;

    #10 $display("\n1 * 2**-51:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3CC0000000000000;

    #10 $display("\n1 * 2**-52:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3CB0000000000000;

    #10 $display("\n1 * 2**-53:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3CA0000000000000;

    #10 $display("\n1 * 2**-54:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3C90000000000000;

    #10 $display("\n1 * 2**-55:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3C80000000000000;

    #10 $display("\n1 * 2**-56:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3C70000000000000;

    #10 $display("\n1 * 2**-57:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3C60000000000000;

    #10 $display("\n1 * 2**-58:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3C50000000000000;

    #10 $display("\n1 * 2**-59:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3C40000000000000;

    #10 $display("\n1 * 2**-60:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3C30000000000000;

    #10 $display("\n1 * 2**-61:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3C20000000000000;

    #10 $display("\n1 * 2**-62:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3C10000000000000;

    #10 $display("\n1 * 2**-63:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3C00000000000000;

    #10 $display("\n1 * 2**-64:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3BF0000000000000;

    #10 $display("\n1 * 2**-65:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3BE0000000000000;

    #10 $display("\n1 * 2**-66:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3BD0000000000000;

    #10 $display("\n1 * 2**-67:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3BC0000000000000;

    #10 $display("\n1 * 2**-68:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3BB0000000000000;

    #10 $display("\n1 * 2**-69:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3BA0000000000000;

    #10 $display("\n1 * 2**-70:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3B90000000000000;

    #10 $display("\n1 * 2**-71:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3B80000000000000;

    #10 $display("\n1 * 2**-72:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3B70000000000000;

    #10 $display("\n1 * 2**-73:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3B60000000000000;

    #10 $display("\n1 * 2**-74:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3B50000000000000;

    #10 $display("\n1 * 2**-75:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3B40000000000000;

    #10 $display("\n1 * 2**-76:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3B30000000000000;

    #10 $display("\n1 * 2**-77:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3B20000000000000;

    #10 $display("\n1 * 2**-78:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3B10000000000000;

    #10 $display("\n1 * 2**-79:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3B00000000000000;

    #10 $display("\n1 * 2**-80:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3AF0000000000000;

    #10 $display("\n1 * 2**-81:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3AE0000000000000;

    #10 $display("\n1 * 2**-82:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3AD0000000000000;

    #10 $display("\n1 * 2**-83:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3AC0000000000000;

    #10 $display("\n1 * 2**-84:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3AB0000000000000;

    #10 $display("\n1 * 2**-85:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3AA0000000000000;

    #10 $display("\n1 * 2**-86:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3A90000000000000;

    #10 $display("\n1 * 2**-87:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3A80000000000000;

    #10 $display("\n1 * 2**-88:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3A70000000000000;

    #10 $display("\n1 * 2**-89:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3A60000000000000;

    #10 $display("\n1 * 2**-90:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3A50000000000000;

    #10 $display("\n1 * 2**-91:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3A40000000000000;

    #10 $display("\n1 * 2**-92:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3A30000000000000;

    #10 $display("\n1 * 2**-93:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3A20000000000000;

    #10 $display("\n1 * 2**-94:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3A10000000000000;

    #10 $display("\n1 * 2**-95:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3A00000000000000;

    #10 $display("\n1 * 2**-96:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h39F0000000000000;

    #10 $display("\n1 * 2**-97:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h39E0000000000000;

    #10 $display("\n1 * 2**-98:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h39D0000000000000;

    #10 $display("\n1 * 2**-99:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h39C0000000000000;

    #10 $display("\n1 * 2**-100:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h39B0000000000000;

    #10 $display("\n1 * 2**-101:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h39A0000000000000;

    #10 $display("\n1 * 2**-102:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3990000000000000;

    #10 $display("\n1 * 2**-103:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3980000000000000;

    #10 $display("\n1 * 2**-104:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3970000000000000;

    #10 $display("\n1 * 2**-105:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3960000000000000;

    #10 $display("\n1 * 2**-106:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3950000000000000;

    #10 $display("\n1 * 2**-107:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3940000000000000;

    #10 $display("\n1 * 2**-108:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3930000000000000;

    #10 $display("\n1 * 2**-109:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3920000000000000;

    #10 $display("\n1 * 2**-110:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3910000000000000;

    #10 $display("\n1 * 2**-111:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3900000000000000;

    #10 $display("\n1 * 2**-112:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h38F0000000000000;

    #10 $display("\n1 * 2**-113:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h38E0000000000000;

    #10 $display("\n1 * 2**-114:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h38D0000000000000;

    #10 $display("\n1 * 2**-115:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h38C0000000000000;

    #10 $display("\n1 * 2**-116:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h38B0000000000000;

    #10 $display("\n1 * 2**-117:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h38A0000000000000;

    #10 $display("\n1 * 2**-118:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3890000000000000;

    #10 $display("\n1 * 2**-119:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3880000000000000;

    #10 $display("\n1 * 2**-120:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3870000000000000;

    #10 $display("\n1 * 2**-121:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3860000000000000;

    #10 $display("\n1 * 2**-122:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3850000000000000;

    #10 $display("\n1 * 2**-123:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3840000000000000;

    #10 $display("\n1 * 2**-124:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3830000000000000;

    #10 $display("\n1 * 2**-125:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3820000000000000;

    #10 $display("\n1 * 2**-126:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3810000000000000;

    #10 $display("\n1 * 2**-127:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3800000000000000;

    #10 $display("\n1 * 2**-128:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h37F0000000000000;

    #10 $display("\n1 * 2**-129:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h37E0000000000000;

    #10 $display("\n1 * 2**-130:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h37D0000000000000;

    #10 $display("\n1 * 2**-131:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h37C0000000000000;

    #10 $display("\n1 * 2**-132:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h37B0000000000000;

    #10 $display("\n1 * 2**-133:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h37A0000000000000;

    #10 $display("\n1 * 2**-134:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3790000000000000;

    #10 $display("\n1 * 2**-135:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3780000000000000;

    #10 $display("\n1 * 2**-136:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3770000000000000;

    #10 $display("\n1 * 2**-137:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3760000000000000;

    #10 $display("\n1 * 2**-138:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3750000000000000;

    #10 $display("\n1 * 2**-139:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3740000000000000;

    #10 $display("\n1 * 2**-140:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3730000000000000;

    #10 $display("\n1 * 2**-141:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3720000000000000;

    #10 $display("\n1 * 2**-142:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3710000000000000;

    #10 $display("\n1 * 2**-143:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3700000000000000;

    #10 $display("\n1 * 2**-144:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h36F0000000000000;

    #10 $display("\n1 * 2**-145:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h36E0000000000000;

    #10 $display("\n1 * 2**-146:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h36D0000000000000;

    #10 $display("\n1 * 2**-147:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h36C0000000000000;

    #10 $display("\n1 * 2**-148:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h36B0000000000000;

    #10 $display("\n1 * 2**-149:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h36A0000000000000;

    #10 $display("\n1 * 2**-150:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3690000000000000;

    #10 $display("\n1 * 2**-151:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3680000000000000;

    #10 $display("\n1 * 2**-152:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3670000000000000;

    #10 $display("\n1 * 2**-153:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3660000000000000;

    #10 $display("\n1 * 2**-154:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3650000000000000;

    #10 $display("\n1 * 2**-155:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3640000000000000;

    #10 $display("\n1 * 2**-156:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3630000000000000;

    #10 $display("\n1 * 2**-157:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3620000000000000;

    #10 $display("\n1 * 2**-158:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3610000000000000;

    #10 $display("\n1 * 2**-159:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3600000000000000;

    #10 $display("\n1 * 2**-160:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h35F0000000000000;

    #10 $display("\n1 * 2**-161:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h35E0000000000000;

    #10 $display("\n1 * 2**-162:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h35D0000000000000;

    #10 $display("\n1 * 2**-163:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h35C0000000000000;

    #10 $display("\n1 * 2**-164:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h35B0000000000000;

    #10 $display("\n1 * 2**-165:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h35A0000000000000;

    #10 $display("\n1 * 2**-166:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3590000000000000;

    #10 $display("\n1 * 2**-167:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3580000000000000;

    #10 $display("\n1 * 2**-168:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3570000000000000;

    #10 $display("\n1 * 2**-169:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3560000000000000;

    #10 $display("\n1 * 2**-170:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3550000000000000;

    #10 $display("\n1 * 2**-171:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3540000000000000;

    #10 $display("\n1 * 2**-172:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3530000000000000;

    #10 $display("\n1 * 2**-173:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3520000000000000;

    #10 $display("\n1 * 2**-174:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3510000000000000;

    #10 $display("\n1 * 2**-175:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3500000000000000;

    #10 $display("\n1 * 2**-176:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h34F0000000000000;

    #10 $display("\n1 * 2**-177:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h34E0000000000000;

    #10 $display("\n1 * 2**-178:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h34D0000000000000;

    #10 $display("\n1 * 2**-179:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h34C0000000000000;

    #10 $display("\n1 * 2**-180:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h34B0000000000000;

    #10 $display("\n1 * 2**-181:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h34A0000000000000;

    #10 $display("\n1 * 2**-182:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3490000000000000;

    #10 $display("\n1 * 2**-183:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3480000000000000;

    #10 $display("\n1 * 2**-184:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3470000000000000;

    #10 $display("\n1 * 2**-185:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3460000000000000;

    #10 $display("\n1 * 2**-186:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3450000000000000;

    #10 $display("\n1 * 2**-187:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3440000000000000;

    #10 $display("\n1 * 2**-188:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3430000000000000;

    #10 $display("\n1 * 2**-189:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3420000000000000;

    #10 $display("\n1 * 2**-190:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3410000000000000;

    #10 $display("\n1 * 2**-191:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3400000000000000;

    #10 $display("\n1 * 2**-192:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h33F0000000000000;

    #10 $display("\n1 * 2**-193:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h33E0000000000000;

    #10 $display("\n1 * 2**-194:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h33D0000000000000;

    #10 $display("\n1 * 2**-195:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h33C0000000000000;

    #10 $display("\n1 * 2**-196:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h33B0000000000000;

    #10 $display("\n1 * 2**-197:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h33A0000000000000;

    #10 $display("\n1 * 2**-198:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3390000000000000;

    #10 $display("\n1 * 2**-199:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3380000000000000;

    #10 $display("\n1 * 2**-200:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3370000000000000;

    #10 $display("\n1 * 2**-201:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3360000000000000;

    #10 $display("\n1 * 2**-202:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3350000000000000;

    #10 $display("\n1 * 2**-203:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3340000000000000;

    #10 $display("\n1 * 2**-204:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3330000000000000;

    #10 $display("\n1 * 2**-205:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3320000000000000;

    #10 $display("\n1 * 2**-206:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3310000000000000;

    #10 $display("\n1 * 2**-207:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3300000000000000;

    #10 $display("\n1 * 2**-208:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h32F0000000000000;

    #10 $display("\n1 * 2**-209:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h32E0000000000000;

    #10 $display("\n1 * 2**-210:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h32D0000000000000;

    #10 $display("\n1 * 2**-211:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h32C0000000000000;

    #10 $display("\n1 * 2**-212:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h32B0000000000000;

    #10 $display("\n1 * 2**-213:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h32A0000000000000;

    #10 $display("\n1 * 2**-214:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3290000000000000;

    #10 $display("\n1 * 2**-215:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3280000000000000;

    #10 $display("\n1 * 2**-216:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3270000000000000;

    #10 $display("\n1 * 2**-217:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3260000000000000;

    #10 $display("\n1 * 2**-218:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3250000000000000;

    #10 $display("\n1 * 2**-219:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3240000000000000;

    #10 $display("\n1 * 2**-220:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3230000000000000;

    #10 $display("\n1 * 2**-221:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3220000000000000;

    #10 $display("\n1 * 2**-222:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3210000000000000;

    #10 $display("\n1 * 2**-223:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3200000000000000;

    #10 $display("\n1 * 2**-224:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h31F0000000000000;

    #10 $display("\n1 * 2**-225:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h31E0000000000000;

    #10 $display("\n1 * 2**-226:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h31D0000000000000;

    #10 $display("\n1 * 2**-227:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h31C0000000000000;

    #10 $display("\n1 * 2**-228:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h31B0000000000000;

    #10 $display("\n1 * 2**-229:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h31A0000000000000;

    #10 $display("\n1 * 2**-230:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3190000000000000;

    #10 $display("\n1 * 2**-231:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3180000000000000;

    #10 $display("\n1 * 2**-232:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3170000000000000;

    #10 $display("\n1 * 2**-233:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3160000000000000;

    #10 $display("\n1 * 2**-234:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3150000000000000;

    #10 $display("\n1 * 2**-235:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3140000000000000;

    #10 $display("\n1 * 2**-236:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3130000000000000;

    #10 $display("\n1 * 2**-237:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3120000000000000;

    #10 $display("\n1 * 2**-238:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3110000000000000;

    #10 $display("\n1 * 2**-239:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3100000000000000;

    #10 $display("\n1 * 2**-240:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h30F0000000000000;

    #10 $display("\n1 * 2**-241:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h30E0000000000000;

    #10 $display("\n1 * 2**-242:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h30D0000000000000;

    #10 $display("\n1 * 2**-243:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h30C0000000000000;

    #10 $display("\n1 * 2**-244:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h30B0000000000000;

    #10 $display("\n1 * 2**-245:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h30A0000000000000;

    #10 $display("\n1 * 2**-246:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3090000000000000;

    #10 $display("\n1 * 2**-247:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3080000000000000;

    #10 $display("\n1 * 2**-248:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3070000000000000;

    #10 $display("\n1 * 2**-249:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3060000000000000;

    #10 $display("\n1 * 2**-250:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3050000000000000;

    #10 $display("\n1 * 2**-251:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3040000000000000;

    #10 $display("\n1 * 2**-252:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3030000000000000;

    #10 $display("\n1 * 2**-253:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3020000000000000;

    #10 $display("\n1 * 2**-254:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3010000000000000;

    #10 $display("\n1 * 2**-255:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h3000000000000000;

    #10 $display("\n1 * 2**-256:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2FF0000000000000;

    #10 $display("\n1 * 2**-257:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2FE0000000000000;

    #10 $display("\n1 * 2**-258:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2FD0000000000000;

    #10 $display("\n1 * 2**-259:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2FC0000000000000;

    #10 $display("\n1 * 2**-260:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2FB0000000000000;

    #10 $display("\n1 * 2**-261:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2FA0000000000000;

    #10 $display("\n1 * 2**-262:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2F90000000000000;

    #10 $display("\n1 * 2**-263:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2F80000000000000;

    #10 $display("\n1 * 2**-264:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2F70000000000000;

    #10 $display("\n1 * 2**-265:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2F60000000000000;

    #10 $display("\n1 * 2**-266:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2F50000000000000;

    #10 $display("\n1 * 2**-267:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2F40000000000000;

    #10 $display("\n1 * 2**-268:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2F30000000000000;

    #10 $display("\n1 * 2**-269:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2F20000000000000;

    #10 $display("\n1 * 2**-270:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2F10000000000000;

    #10 $display("\n1 * 2**-271:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2F00000000000000;

    #10 $display("\n1 * 2**-272:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2EF0000000000000;

    #10 $display("\n1 * 2**-273:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2EE0000000000000;

    #10 $display("\n1 * 2**-274:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2ED0000000000000;

    #10 $display("\n1 * 2**-275:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2EC0000000000000;

    #10 $display("\n1 * 2**-276:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2EB0000000000000;

    #10 $display("\n1 * 2**-277:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2EA0000000000000;

    #10 $display("\n1 * 2**-278:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2E90000000000000;

    #10 $display("\n1 * 2**-279:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2E80000000000000;

    #10 $display("\n1 * 2**-280:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2E70000000000000;

    #10 $display("\n1 * 2**-281:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2E60000000000000;

    #10 $display("\n1 * 2**-282:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2E50000000000000;

    #10 $display("\n1 * 2**-283:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2E40000000000000;

    #10 $display("\n1 * 2**-284:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2E30000000000000;

    #10 $display("\n1 * 2**-285:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2E20000000000000;

    #10 $display("\n1 * 2**-286:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2E10000000000000;

    #10 $display("\n1 * 2**-287:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2E00000000000000;

    #10 $display("\n1 * 2**-288:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2DF0000000000000;

    #10 $display("\n1 * 2**-289:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2DE0000000000000;

    #10 $display("\n1 * 2**-290:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2DD0000000000000;

    #10 $display("\n1 * 2**-291:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2DC0000000000000;

    #10 $display("\n1 * 2**-292:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2DB0000000000000;

    #10 $display("\n1 * 2**-293:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2DA0000000000000;

    #10 $display("\n1 * 2**-294:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2D90000000000000;

    #10 $display("\n1 * 2**-295:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2D80000000000000;

    #10 $display("\n1 * 2**-296:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2D70000000000000;

    #10 $display("\n1 * 2**-297:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2D60000000000000;

    #10 $display("\n1 * 2**-298:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2D50000000000000;

    #10 $display("\n1 * 2**-299:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2D40000000000000;

    #10 $display("\n1 * 2**-300:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2D30000000000000;

    #10 $display("\n1 * 2**-301:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2D20000000000000;

    #10 $display("\n1 * 2**-302:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2D10000000000000;

    #10 $display("\n1 * 2**-303:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2D00000000000000;

    #10 $display("\n1 * 2**-304:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2CF0000000000000;

    #10 $display("\n1 * 2**-305:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2CE0000000000000;

    #10 $display("\n1 * 2**-306:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2CD0000000000000;

    #10 $display("\n1 * 2**-307:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2CC0000000000000;

    #10 $display("\n1 * 2**-308:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2CB0000000000000;

    #10 $display("\n1 * 2**-309:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2CA0000000000000;

    #10 $display("\n1 * 2**-310:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2C90000000000000;

    #10 $display("\n1 * 2**-311:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2C80000000000000;

    #10 $display("\n1 * 2**-312:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2C70000000000000;

    #10 $display("\n1 * 2**-313:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2C60000000000000;

    #10 $display("\n1 * 2**-314:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2C50000000000000;

    #10 $display("\n1 * 2**-315:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2C40000000000000;

    #10 $display("\n1 * 2**-316:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2C30000000000000;

    #10 $display("\n1 * 2**-317:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2C20000000000000;

    #10 $display("\n1 * 2**-318:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2C10000000000000;

    #10 $display("\n1 * 2**-319:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2C00000000000000;

    #10 $display("\n1 * 2**-320:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2BF0000000000000;

    #10 $display("\n1 * 2**-321:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2BE0000000000000;

    #10 $display("\n1 * 2**-322:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2BD0000000000000;

    #10 $display("\n1 * 2**-323:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2BC0000000000000;

    #10 $display("\n1 * 2**-324:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2BB0000000000000;

    #10 $display("\n1 * 2**-325:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2BA0000000000000;

    #10 $display("\n1 * 2**-326:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2B90000000000000;

    #10 $display("\n1 * 2**-327:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2B80000000000000;

    #10 $display("\n1 * 2**-328:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2B70000000000000;

    #10 $display("\n1 * 2**-329:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2B60000000000000;

    #10 $display("\n1 * 2**-330:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2B50000000000000;

    #10 $display("\n1 * 2**-331:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2B40000000000000;

    #10 $display("\n1 * 2**-332:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2B30000000000000;

    #10 $display("\n1 * 2**-333:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2B20000000000000;

    #10 $display("\n1 * 2**-334:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2B10000000000000;

    #10 $display("\n1 * 2**-335:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2B00000000000000;

    #10 $display("\n1 * 2**-336:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2AF0000000000000;

    #10 $display("\n1 * 2**-337:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2AE0000000000000;

    #10 $display("\n1 * 2**-338:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2AD0000000000000;

    #10 $display("\n1 * 2**-339:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2AC0000000000000;

    #10 $display("\n1 * 2**-340:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2AB0000000000000;

    #10 $display("\n1 * 2**-341:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2AA0000000000000;

    #10 $display("\n1 * 2**-342:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2A90000000000000;

    #10 $display("\n1 * 2**-343:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2A80000000000000;

    #10 $display("\n1 * 2**-344:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2A70000000000000;

    #10 $display("\n1 * 2**-345:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2A60000000000000;

    #10 $display("\n1 * 2**-346:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2A50000000000000;

    #10 $display("\n1 * 2**-347:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2A40000000000000;

    #10 $display("\n1 * 2**-348:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2A30000000000000;

    #10 $display("\n1 * 2**-349:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2A20000000000000;

    #10 $display("\n1 * 2**-350:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2A10000000000000;

    #10 $display("\n1 * 2**-351:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2A00000000000000;

    #10 $display("\n1 * 2**-352:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h29F0000000000000;

    #10 $display("\n1 * 2**-353:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h29E0000000000000;

    #10 $display("\n1 * 2**-354:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h29D0000000000000;

    #10 $display("\n1 * 2**-355:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h29C0000000000000;

    #10 $display("\n1 * 2**-356:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h29B0000000000000;

    #10 $display("\n1 * 2**-357:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h29A0000000000000;

    #10 $display("\n1 * 2**-358:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2990000000000000;

    #10 $display("\n1 * 2**-359:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2980000000000000;

    #10 $display("\n1 * 2**-360:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2970000000000000;

    #10 $display("\n1 * 2**-361:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2960000000000000;

    #10 $display("\n1 * 2**-362:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2950000000000000;

    #10 $display("\n1 * 2**-363:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2940000000000000;

    #10 $display("\n1 * 2**-364:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2930000000000000;

    #10 $display("\n1 * 2**-365:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2920000000000000;

    #10 $display("\n1 * 2**-366:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2910000000000000;

    #10 $display("\n1 * 2**-367:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2900000000000000;

    #10 $display("\n1 * 2**-368:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h28F0000000000000;

    #10 $display("\n1 * 2**-369:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h28E0000000000000;

    #10 $display("\n1 * 2**-370:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h28D0000000000000;

    #10 $display("\n1 * 2**-371:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h28C0000000000000;

    #10 $display("\n1 * 2**-372:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h28B0000000000000;

    #10 $display("\n1 * 2**-373:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h28A0000000000000;

    #10 $display("\n1 * 2**-374:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2890000000000000;

    #10 $display("\n1 * 2**-375:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2880000000000000;

    #10 $display("\n1 * 2**-376:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2870000000000000;

    #10 $display("\n1 * 2**-377:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2860000000000000;

    #10 $display("\n1 * 2**-378:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2850000000000000;

    #10 $display("\n1 * 2**-379:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2840000000000000;

    #10 $display("\n1 * 2**-380:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2830000000000000;

    #10 $display("\n1 * 2**-381:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2820000000000000;

    #10 $display("\n1 * 2**-382:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2810000000000000;

    #10 $display("\n1 * 2**-383:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2800000000000000;

    #10 $display("\n1 * 2**-384:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h27F0000000000000;

    #10 $display("\n1 * 2**-385:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h27E0000000000000;

    #10 $display("\n1 * 2**-386:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h27D0000000000000;

    #10 $display("\n1 * 2**-387:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h27C0000000000000;

    #10 $display("\n1 * 2**-388:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h27B0000000000000;

    #10 $display("\n1 * 2**-389:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h27A0000000000000;

    #10 $display("\n1 * 2**-390:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2790000000000000;

    #10 $display("\n1 * 2**-391:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2780000000000000;

    #10 $display("\n1 * 2**-392:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2770000000000000;

    #10 $display("\n1 * 2**-393:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2760000000000000;

    #10 $display("\n1 * 2**-394:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2750000000000000;

    #10 $display("\n1 * 2**-395:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2740000000000000;

    #10 $display("\n1 * 2**-396:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2730000000000000;

    #10 $display("\n1 * 2**-397:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2720000000000000;

    #10 $display("\n1 * 2**-398:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2710000000000000;

    #10 $display("\n1 * 2**-399:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2700000000000000;

    #10 $display("\n1 * 2**-400:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h26F0000000000000;

    #10 $display("\n1 * 2**-401:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h26E0000000000000;

    #10 $display("\n1 * 2**-402:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h26D0000000000000;

    #10 $display("\n1 * 2**-403:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h26C0000000000000;

    #10 $display("\n1 * 2**-404:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h26B0000000000000;

    #10 $display("\n1 * 2**-405:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h26A0000000000000;

    #10 $display("\n1 * 2**-406:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2690000000000000;

    #10 $display("\n1 * 2**-407:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2680000000000000;

    #10 $display("\n1 * 2**-408:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2670000000000000;

    #10 $display("\n1 * 2**-409:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2660000000000000;

    #10 $display("\n1 * 2**-410:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2650000000000000;

    #10 $display("\n1 * 2**-411:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2640000000000000;

    #10 $display("\n1 * 2**-412:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2630000000000000;

    #10 $display("\n1 * 2**-413:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2620000000000000;

    #10 $display("\n1 * 2**-414:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2610000000000000;

    #10 $display("\n1 * 2**-415:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2600000000000000;

    #10 $display("\n1 * 2**-416:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h25F0000000000000;

    #10 $display("\n1 * 2**-417:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h25E0000000000000;

    #10 $display("\n1 * 2**-418:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h25D0000000000000;

    #10 $display("\n1 * 2**-419:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h25C0000000000000;

    #10 $display("\n1 * 2**-420:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h25B0000000000000;

    #10 $display("\n1 * 2**-421:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h25A0000000000000;

    #10 $display("\n1 * 2**-422:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2590000000000000;

    #10 $display("\n1 * 2**-423:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2580000000000000;

    #10 $display("\n1 * 2**-424:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2570000000000000;

    #10 $display("\n1 * 2**-425:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2560000000000000;

    #10 $display("\n1 * 2**-426:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2550000000000000;

    #10 $display("\n1 * 2**-427:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2540000000000000;

    #10 $display("\n1 * 2**-428:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2530000000000000;

    #10 $display("\n1 * 2**-429:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2520000000000000;

    #10 $display("\n1 * 2**-430:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2510000000000000;

    #10 $display("\n1 * 2**-431:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2500000000000000;

    #10 $display("\n1 * 2**-432:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h24F0000000000000;

    #10 $display("\n1 * 2**-433:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h24E0000000000000;

    #10 $display("\n1 * 2**-434:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h24D0000000000000;

    #10 $display("\n1 * 2**-435:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h24C0000000000000;

    #10 $display("\n1 * 2**-436:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h24B0000000000000;

    #10 $display("\n1 * 2**-437:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h24A0000000000000;

    #10 $display("\n1 * 2**-438:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2490000000000000;

    #10 $display("\n1 * 2**-439:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2480000000000000;

    #10 $display("\n1 * 2**-440:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2470000000000000;

    #10 $display("\n1 * 2**-441:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2460000000000000;

    #10 $display("\n1 * 2**-442:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2450000000000000;

    #10 $display("\n1 * 2**-443:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2440000000000000;

    #10 $display("\n1 * 2**-444:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2430000000000000;

    #10 $display("\n1 * 2**-445:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2420000000000000;

    #10 $display("\n1 * 2**-446:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2410000000000000;

    #10 $display("\n1 * 2**-447:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2400000000000000;

    #10 $display("\n1 * 2**-448:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h23F0000000000000;

    #10 $display("\n1 * 2**-449:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h23E0000000000000;

    #10 $display("\n1 * 2**-450:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h23D0000000000000;

    #10 $display("\n1 * 2**-451:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h23C0000000000000;

    #10 $display("\n1 * 2**-452:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h23B0000000000000;

    #10 $display("\n1 * 2**-453:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h23A0000000000000;

    #10 $display("\n1 * 2**-454:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2390000000000000;

    #10 $display("\n1 * 2**-455:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2380000000000000;

    #10 $display("\n1 * 2**-456:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2370000000000000;

    #10 $display("\n1 * 2**-457:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2360000000000000;

    #10 $display("\n1 * 2**-458:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2350000000000000;

    #10 $display("\n1 * 2**-459:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2340000000000000;

    #10 $display("\n1 * 2**-460:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2330000000000000;

    #10 $display("\n1 * 2**-461:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2320000000000000;

    #10 $display("\n1 * 2**-462:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2310000000000000;

    #10 $display("\n1 * 2**-463:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2300000000000000;

    #10 $display("\n1 * 2**-464:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h22F0000000000000;

    #10 $display("\n1 * 2**-465:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h22E0000000000000;

    #10 $display("\n1 * 2**-466:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h22D0000000000000;

    #10 $display("\n1 * 2**-467:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h22C0000000000000;

    #10 $display("\n1 * 2**-468:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h22B0000000000000;

    #10 $display("\n1 * 2**-469:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h22A0000000000000;

    #10 $display("\n1 * 2**-470:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2290000000000000;

    #10 $display("\n1 * 2**-471:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2280000000000000;

    #10 $display("\n1 * 2**-472:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2270000000000000;

    #10 $display("\n1 * 2**-473:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2260000000000000;

    #10 $display("\n1 * 2**-474:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2250000000000000;

    #10 $display("\n1 * 2**-475:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2240000000000000;

    #10 $display("\n1 * 2**-476:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2230000000000000;

    #10 $display("\n1 * 2**-477:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2220000000000000;

    #10 $display("\n1 * 2**-478:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2210000000000000;

    #10 $display("\n1 * 2**-479:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2200000000000000;

    #10 $display("\n1 * 2**-480:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h21F0000000000000;

    #10 $display("\n1 * 2**-481:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h21E0000000000000;

    #10 $display("\n1 * 2**-482:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h21D0000000000000;

    #10 $display("\n1 * 2**-483:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h21C0000000000000;

    #10 $display("\n1 * 2**-484:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h21B0000000000000;

    #10 $display("\n1 * 2**-485:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h21A0000000000000;

    #10 $display("\n1 * 2**-486:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2190000000000000;

    #10 $display("\n1 * 2**-487:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2180000000000000;

    #10 $display("\n1 * 2**-488:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2170000000000000;

    #10 $display("\n1 * 2**-489:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2160000000000000;

    #10 $display("\n1 * 2**-490:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2150000000000000;

    #10 $display("\n1 * 2**-491:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2140000000000000;

    #10 $display("\n1 * 2**-492:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2130000000000000;

    #10 $display("\n1 * 2**-493:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2120000000000000;

    #10 $display("\n1 * 2**-494:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2110000000000000;

    #10 $display("\n1 * 2**-495:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2100000000000000;

    #10 $display("\n1 * 2**-496:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h20F0000000000000;

    #10 $display("\n1 * 2**-497:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h20E0000000000000;

    #10 $display("\n1 * 2**-498:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h20D0000000000000;

    #10 $display("\n1 * 2**-499:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h20C0000000000000;

    #10 $display("\n1 * 2**-500:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h20B0000000000000;

    #10 $display("\n1 * 2**-501:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h20A0000000000000;

    #10 $display("\n1 * 2**-502:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2090000000000000;

    #10 $display("\n1 * 2**-503:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2080000000000000;

    #10 $display("\n1 * 2**-504:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2070000000000000;

    #10 $display("\n1 * 2**-505:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2060000000000000;

    #10 $display("\n1 * 2**-506:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2050000000000000;

    #10 $display("\n1 * 2**-507:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2040000000000000;

    #10 $display("\n1 * 2**-508:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2030000000000000;

    #10 $display("\n1 * 2**-509:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2020000000000000;

    #10 $display("\n1 * 2**-510:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2010000000000000;

    #10 $display("\n1 * 2**-511:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h2000000000000000;

    #10 $display("\n1 * 2**-512:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1FF0000000000000;

    #10 $display("\n1 * 2**-513:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1FE0000000000000;

    #10 $display("\n1 * 2**-514:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1FD0000000000000;

    #10 $display("\n1 * 2**-515:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1FC0000000000000;

    #10 $display("\n1 * 2**-516:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1FB0000000000000;

    #10 $display("\n1 * 2**-517:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1FA0000000000000;

    #10 $display("\n1 * 2**-518:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1F90000000000000;

    #10 $display("\n1 * 2**-519:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1F80000000000000;

    #10 $display("\n1 * 2**-520:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1F70000000000000;

    #10 $display("\n1 * 2**-521:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1F60000000000000;

    #10 $display("\n1 * 2**-522:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1F50000000000000;

    #10 $display("\n1 * 2**-523:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1F40000000000000;

    #10 $display("\n1 * 2**-524:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1F30000000000000;

    #10 $display("\n1 * 2**-525:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1F20000000000000;

    #10 $display("\n1 * 2**-526:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1F10000000000000;

    #10 $display("\n1 * 2**-527:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1F00000000000000;

    #10 $display("\n1 * 2**-528:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1EF0000000000000;

    #10 $display("\n1 * 2**-529:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1EE0000000000000;

    #10 $display("\n1 * 2**-530:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1ED0000000000000;

    #10 $display("\n1 * 2**-531:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1EC0000000000000;

    #10 $display("\n1 * 2**-532:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1EB0000000000000;

    #10 $display("\n1 * 2**-533:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1EA0000000000000;

    #10 $display("\n1 * 2**-534:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1E90000000000000;

    #10 $display("\n1 * 2**-535:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1E80000000000000;

    #10 $display("\n1 * 2**-536:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1E70000000000000;

    #10 $display("\n1 * 2**-537:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1E60000000000000;

    #10 $display("\n1 * 2**-538:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1E50000000000000;

    #10 $display("\n1 * 2**-539:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1E40000000000000;

    #10 $display("\n1 * 2**-540:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1E30000000000000;

    #10 $display("\n1 * 2**-541:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1E20000000000000;

    #10 $display("\n1 * 2**-542:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1E10000000000000;

    #10 $display("\n1 * 2**-543:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1E00000000000000;

    #10 $display("\n1 * 2**-544:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1DF0000000000000;

    #10 $display("\n1 * 2**-545:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1DE0000000000000;

    #10 $display("\n1 * 2**-546:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1DD0000000000000;

    #10 $display("\n1 * 2**-547:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1DC0000000000000;

    #10 $display("\n1 * 2**-548:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1DB0000000000000;

    #10 $display("\n1 * 2**-549:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1DA0000000000000;

    #10 $display("\n1 * 2**-550:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1D90000000000000;

    #10 $display("\n1 * 2**-551:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1D80000000000000;

    #10 $display("\n1 * 2**-552:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1D70000000000000;

    #10 $display("\n1 * 2**-553:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1D60000000000000;

    #10 $display("\n1 * 2**-554:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1D50000000000000;

    #10 $display("\n1 * 2**-555:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1D40000000000000;

    #10 $display("\n1 * 2**-556:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1D30000000000000;

    #10 $display("\n1 * 2**-557:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1D20000000000000;

    #10 $display("\n1 * 2**-558:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1D10000000000000;

    #10 $display("\n1 * 2**-559:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1D00000000000000;

    #10 $display("\n1 * 2**-560:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1CF0000000000000;

    #10 $display("\n1 * 2**-561:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1CE0000000000000;

    #10 $display("\n1 * 2**-562:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1CD0000000000000;

    #10 $display("\n1 * 2**-563:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1CC0000000000000;

    #10 $display("\n1 * 2**-564:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1CB0000000000000;

    #10 $display("\n1 * 2**-565:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1CA0000000000000;

    #10 $display("\n1 * 2**-566:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1C90000000000000;

    #10 $display("\n1 * 2**-567:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1C80000000000000;

    #10 $display("\n1 * 2**-568:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1C70000000000000;

    #10 $display("\n1 * 2**-569:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1C60000000000000;

    #10 $display("\n1 * 2**-570:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1C50000000000000;

    #10 $display("\n1 * 2**-571:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1C40000000000000;

    #10 $display("\n1 * 2**-572:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1C30000000000000;

    #10 $display("\n1 * 2**-573:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1C20000000000000;

    #10 $display("\n1 * 2**-574:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1C10000000000000;

    #10 $display("\n1 * 2**-575:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1C00000000000000;

    #10 $display("\n1 * 2**-576:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1BF0000000000000;

    #10 $display("\n1 * 2**-577:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1BE0000000000000;

    #10 $display("\n1 * 2**-578:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1BD0000000000000;

    #10 $display("\n1 * 2**-579:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1BC0000000000000;

    #10 $display("\n1 * 2**-580:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1BB0000000000000;

    #10 $display("\n1 * 2**-581:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1BA0000000000000;

    #10 $display("\n1 * 2**-582:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1B90000000000000;

    #10 $display("\n1 * 2**-583:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1B80000000000000;

    #10 $display("\n1 * 2**-584:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1B70000000000000;

    #10 $display("\n1 * 2**-585:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1B60000000000000;

    #10 $display("\n1 * 2**-586:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1B50000000000000;

    #10 $display("\n1 * 2**-587:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1B40000000000000;

    #10 $display("\n1 * 2**-588:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1B30000000000000;

    #10 $display("\n1 * 2**-589:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1B20000000000000;

    #10 $display("\n1 * 2**-590:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1B10000000000000;

    #10 $display("\n1 * 2**-591:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1B00000000000000;

    #10 $display("\n1 * 2**-592:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1AF0000000000000;

    #10 $display("\n1 * 2**-593:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1AE0000000000000;

    #10 $display("\n1 * 2**-594:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1AD0000000000000;

    #10 $display("\n1 * 2**-595:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1AC0000000000000;

    #10 $display("\n1 * 2**-596:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1AB0000000000000;

    #10 $display("\n1 * 2**-597:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1AA0000000000000;

    #10 $display("\n1 * 2**-598:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1A90000000000000;

    #10 $display("\n1 * 2**-599:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1A80000000000000;

    #10 $display("\n1 * 2**-600:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1A70000000000000;

    #10 $display("\n1 * 2**-601:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1A60000000000000;

    #10 $display("\n1 * 2**-602:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1A50000000000000;

    #10 $display("\n1 * 2**-603:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1A40000000000000;

    #10 $display("\n1 * 2**-604:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1A30000000000000;

    #10 $display("\n1 * 2**-605:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1A20000000000000;

    #10 $display("\n1 * 2**-606:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1A10000000000000;

    #10 $display("\n1 * 2**-607:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1A00000000000000;

    #10 $display("\n1 * 2**-608:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h19F0000000000000;

    #10 $display("\n1 * 2**-609:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h19E0000000000000;

    #10 $display("\n1 * 2**-610:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h19D0000000000000;

    #10 $display("\n1 * 2**-611:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h19C0000000000000;

    #10 $display("\n1 * 2**-612:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h19B0000000000000;

    #10 $display("\n1 * 2**-613:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h19A0000000000000;

    #10 $display("\n1 * 2**-614:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1990000000000000;

    #10 $display("\n1 * 2**-615:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1980000000000000;

    #10 $display("\n1 * 2**-616:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1970000000000000;

    #10 $display("\n1 * 2**-617:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1960000000000000;

    #10 $display("\n1 * 2**-618:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1950000000000000;

    #10 $display("\n1 * 2**-619:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1940000000000000;

    #10 $display("\n1 * 2**-620:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1930000000000000;

    #10 $display("\n1 * 2**-621:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1920000000000000;

    #10 $display("\n1 * 2**-622:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1910000000000000;

    #10 $display("\n1 * 2**-623:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1900000000000000;

    #10 $display("\n1 * 2**-624:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h18F0000000000000;

    #10 $display("\n1 * 2**-625:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h18E0000000000000;

    #10 $display("\n1 * 2**-626:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h18D0000000000000;

    #10 $display("\n1 * 2**-627:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h18C0000000000000;

    #10 $display("\n1 * 2**-628:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h18B0000000000000;

    #10 $display("\n1 * 2**-629:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h18A0000000000000;

    #10 $display("\n1 * 2**-630:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1890000000000000;

    #10 $display("\n1 * 2**-631:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1880000000000000;

    #10 $display("\n1 * 2**-632:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1870000000000000;

    #10 $display("\n1 * 2**-633:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1860000000000000;

    #10 $display("\n1 * 2**-634:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1850000000000000;

    #10 $display("\n1 * 2**-635:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1840000000000000;

    #10 $display("\n1 * 2**-636:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1830000000000000;

    #10 $display("\n1 * 2**-637:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1820000000000000;

    #10 $display("\n1 * 2**-638:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1810000000000000;

    #10 $display("\n1 * 2**-639:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1800000000000000;

    #10 $display("\n1 * 2**-640:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h17F0000000000000;

    #10 $display("\n1 * 2**-641:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h17E0000000000000;

    #10 $display("\n1 * 2**-642:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h17D0000000000000;

    #10 $display("\n1 * 2**-643:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h17C0000000000000;

    #10 $display("\n1 * 2**-644:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h17B0000000000000;

    #10 $display("\n1 * 2**-645:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h17A0000000000000;

    #10 $display("\n1 * 2**-646:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1790000000000000;

    #10 $display("\n1 * 2**-647:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1780000000000000;

    #10 $display("\n1 * 2**-648:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1770000000000000;

    #10 $display("\n1 * 2**-649:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1760000000000000;

    #10 $display("\n1 * 2**-650:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1750000000000000;

    #10 $display("\n1 * 2**-651:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1740000000000000;

    #10 $display("\n1 * 2**-652:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1730000000000000;

    #10 $display("\n1 * 2**-653:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1720000000000000;

    #10 $display("\n1 * 2**-654:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1710000000000000;

    #10 $display("\n1 * 2**-655:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1700000000000000;

    #10 $display("\n1 * 2**-656:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h16F0000000000000;

    #10 $display("\n1 * 2**-657:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h16E0000000000000;

    #10 $display("\n1 * 2**-658:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h16D0000000000000;

    #10 $display("\n1 * 2**-659:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h16C0000000000000;

    #10 $display("\n1 * 2**-660:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h16B0000000000000;

    #10 $display("\n1 * 2**-661:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h16A0000000000000;

    #10 $display("\n1 * 2**-662:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1690000000000000;

    #10 $display("\n1 * 2**-663:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1680000000000000;

    #10 $display("\n1 * 2**-664:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1670000000000000;

    #10 $display("\n1 * 2**-665:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1660000000000000;

    #10 $display("\n1 * 2**-666:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1650000000000000;

    #10 $display("\n1 * 2**-667:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1640000000000000;

    #10 $display("\n1 * 2**-668:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1630000000000000;

    #10 $display("\n1 * 2**-669:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1620000000000000;

    #10 $display("\n1 * 2**-670:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1610000000000000;

    #10 $display("\n1 * 2**-671:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1600000000000000;

    #10 $display("\n1 * 2**-672:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h15F0000000000000;

    #10 $display("\n1 * 2**-673:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h15E0000000000000;

    #10 $display("\n1 * 2**-674:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h15D0000000000000;

    #10 $display("\n1 * 2**-675:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h15C0000000000000;

    #10 $display("\n1 * 2**-676:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h15B0000000000000;

    #10 $display("\n1 * 2**-677:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h15A0000000000000;

    #10 $display("\n1 * 2**-678:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1590000000000000;

    #10 $display("\n1 * 2**-679:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1580000000000000;

    #10 $display("\n1 * 2**-680:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1570000000000000;

    #10 $display("\n1 * 2**-681:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1560000000000000;

    #10 $display("\n1 * 2**-682:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1550000000000000;

    #10 $display("\n1 * 2**-683:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1540000000000000;

    #10 $display("\n1 * 2**-684:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1530000000000000;

    #10 $display("\n1 * 2**-685:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1520000000000000;

    #10 $display("\n1 * 2**-686:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1510000000000000;

    #10 $display("\n1 * 2**-687:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1500000000000000;

    #10 $display("\n1 * 2**-688:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h14F0000000000000;

    #10 $display("\n1 * 2**-689:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h14E0000000000000;

    #10 $display("\n1 * 2**-690:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h14D0000000000000;

    #10 $display("\n1 * 2**-691:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h14C0000000000000;

    #10 $display("\n1 * 2**-692:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h14B0000000000000;

    #10 $display("\n1 * 2**-693:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h14A0000000000000;

    #10 $display("\n1 * 2**-694:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1490000000000000;

    #10 $display("\n1 * 2**-695:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1480000000000000;

    #10 $display("\n1 * 2**-696:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1470000000000000;

    #10 $display("\n1 * 2**-697:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1460000000000000;

    #10 $display("\n1 * 2**-698:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1450000000000000;

    #10 $display("\n1 * 2**-699:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1440000000000000;

    #10 $display("\n1 * 2**-700:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1430000000000000;

    #10 $display("\n1 * 2**-701:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1420000000000000;

    #10 $display("\n1 * 2**-702:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1410000000000000;

    #10 $display("\n1 * 2**-703:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1400000000000000;

    #10 $display("\n1 * 2**-704:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h13F0000000000000;

    #10 $display("\n1 * 2**-705:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h13E0000000000000;

    #10 $display("\n1 * 2**-706:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h13D0000000000000;

    #10 $display("\n1 * 2**-707:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h13C0000000000000;

    #10 $display("\n1 * 2**-708:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h13B0000000000000;

    #10 $display("\n1 * 2**-709:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h13A0000000000000;

    #10 $display("\n1 * 2**-710:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1390000000000000;

    #10 $display("\n1 * 2**-711:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1380000000000000;

    #10 $display("\n1 * 2**-712:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1370000000000000;

    #10 $display("\n1 * 2**-713:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1360000000000000;

    #10 $display("\n1 * 2**-714:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1350000000000000;

    #10 $display("\n1 * 2**-715:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1340000000000000;

    #10 $display("\n1 * 2**-716:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1330000000000000;

    #10 $display("\n1 * 2**-717:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1320000000000000;

    #10 $display("\n1 * 2**-718:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1310000000000000;

    #10 $display("\n1 * 2**-719:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1300000000000000;

    #10 $display("\n1 * 2**-720:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h12F0000000000000;

    #10 $display("\n1 * 2**-721:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h12E0000000000000;

    #10 $display("\n1 * 2**-722:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h12D0000000000000;

    #10 $display("\n1 * 2**-723:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h12C0000000000000;

    #10 $display("\n1 * 2**-724:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h12B0000000000000;

    #10 $display("\n1 * 2**-725:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h12A0000000000000;

    #10 $display("\n1 * 2**-726:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1290000000000000;

    #10 $display("\n1 * 2**-727:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1280000000000000;

    #10 $display("\n1 * 2**-728:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1270000000000000;

    #10 $display("\n1 * 2**-729:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1260000000000000;

    #10 $display("\n1 * 2**-730:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1250000000000000;

    #10 $display("\n1 * 2**-731:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1240000000000000;

    #10 $display("\n1 * 2**-732:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1230000000000000;

    #10 $display("\n1 * 2**-733:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1220000000000000;

    #10 $display("\n1 * 2**-734:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1210000000000000;

    #10 $display("\n1 * 2**-735:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1200000000000000;

    #10 $display("\n1 * 2**-736:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h11F0000000000000;

    #10 $display("\n1 * 2**-737:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h11E0000000000000;

    #10 $display("\n1 * 2**-738:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h11D0000000000000;

    #10 $display("\n1 * 2**-739:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h11C0000000000000;

    #10 $display("\n1 * 2**-740:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h11B0000000000000;

    #10 $display("\n1 * 2**-741:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h11A0000000000000;

    #10 $display("\n1 * 2**-742:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1190000000000000;

    #10 $display("\n1 * 2**-743:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1180000000000000;

    #10 $display("\n1 * 2**-744:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1170000000000000;

    #10 $display("\n1 * 2**-745:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1160000000000000;

    #10 $display("\n1 * 2**-746:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1150000000000000;

    #10 $display("\n1 * 2**-747:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1140000000000000;

    #10 $display("\n1 * 2**-748:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1130000000000000;

    #10 $display("\n1 * 2**-749:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1120000000000000;

    #10 $display("\n1 * 2**-750:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1110000000000000;

    #10 $display("\n1 * 2**-751:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1100000000000000;

    #10 $display("\n1 * 2**-752:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h10F0000000000000;

    #10 $display("\n1 * 2**-753:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h10E0000000000000;

    #10 $display("\n1 * 2**-754:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h10D0000000000000;

    #10 $display("\n1 * 2**-755:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h10C0000000000000;

    #10 $display("\n1 * 2**-756:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h10B0000000000000;

    #10 $display("\n1 * 2**-757:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h10A0000000000000;

    #10 $display("\n1 * 2**-758:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1090000000000000;

    #10 $display("\n1 * 2**-759:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1080000000000000;

    #10 $display("\n1 * 2**-760:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1070000000000000;

    #10 $display("\n1 * 2**-761:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1060000000000000;

    #10 $display("\n1 * 2**-762:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1050000000000000;

    #10 $display("\n1 * 2**-763:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1040000000000000;

    #10 $display("\n1 * 2**-764:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1030000000000000;

    #10 $display("\n1 * 2**-765:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1020000000000000;

    #10 $display("\n1 * 2**-766:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1010000000000000;

    #10 $display("\n1 * 2**-767:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h1000000000000000;

    #10 $display("\n1 * 2**-768:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0FF0000000000000;

    #10 $display("\n1 * 2**-769:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0FE0000000000000;

    #10 $display("\n1 * 2**-770:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0FD0000000000000;

    #10 $display("\n1 * 2**-771:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0FC0000000000000;

    #10 $display("\n1 * 2**-772:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0FB0000000000000;

    #10 $display("\n1 * 2**-773:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0FA0000000000000;

    #10 $display("\n1 * 2**-774:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0F90000000000000;

    #10 $display("\n1 * 2**-775:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0F80000000000000;

    #10 $display("\n1 * 2**-776:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0F70000000000000;

    #10 $display("\n1 * 2**-777:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0F60000000000000;

    #10 $display("\n1 * 2**-778:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0F50000000000000;

    #10 $display("\n1 * 2**-779:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0F40000000000000;

    #10 $display("\n1 * 2**-780:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0F30000000000000;

    #10 $display("\n1 * 2**-781:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0F20000000000000;

    #10 $display("\n1 * 2**-782:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0F10000000000000;

    #10 $display("\n1 * 2**-783:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0F00000000000000;

    #10 $display("\n1 * 2**-784:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0EF0000000000000;

    #10 $display("\n1 * 2**-785:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0EE0000000000000;

    #10 $display("\n1 * 2**-786:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0ED0000000000000;

    #10 $display("\n1 * 2**-787:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0EC0000000000000;

    #10 $display("\n1 * 2**-788:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0EB0000000000000;

    #10 $display("\n1 * 2**-789:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0EA0000000000000;

    #10 $display("\n1 * 2**-790:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0E90000000000000;

    #10 $display("\n1 * 2**-791:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0E80000000000000;

    #10 $display("\n1 * 2**-792:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0E70000000000000;

    #10 $display("\n1 * 2**-793:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0E60000000000000;

    #10 $display("\n1 * 2**-794:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0E50000000000000;

    #10 $display("\n1 * 2**-795:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0E40000000000000;

    #10 $display("\n1 * 2**-796:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0E30000000000000;

    #10 $display("\n1 * 2**-797:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0E20000000000000;

    #10 $display("\n1 * 2**-798:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0E10000000000000;

    #10 $display("\n1 * 2**-799:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0E00000000000000;

    #10 $display("\n1 * 2**-800:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0DF0000000000000;

    #10 $display("\n1 * 2**-801:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0DE0000000000000;

    #10 $display("\n1 * 2**-802:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0DD0000000000000;

    #10 $display("\n1 * 2**-803:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0DC0000000000000;

    #10 $display("\n1 * 2**-804:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0DB0000000000000;

    #10 $display("\n1 * 2**-805:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0DA0000000000000;

    #10 $display("\n1 * 2**-806:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0D90000000000000;

    #10 $display("\n1 * 2**-807:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0D80000000000000;

    #10 $display("\n1 * 2**-808:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0D70000000000000;

    #10 $display("\n1 * 2**-809:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0D60000000000000;

    #10 $display("\n1 * 2**-810:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0D50000000000000;

    #10 $display("\n1 * 2**-811:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0D40000000000000;

    #10 $display("\n1 * 2**-812:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0D30000000000000;

    #10 $display("\n1 * 2**-813:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0D20000000000000;

    #10 $display("\n1 * 2**-814:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0D10000000000000;

    #10 $display("\n1 * 2**-815:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0D00000000000000;

    #10 $display("\n1 * 2**-816:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0CF0000000000000;

    #10 $display("\n1 * 2**-817:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0CE0000000000000;

    #10 $display("\n1 * 2**-818:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0CD0000000000000;

    #10 $display("\n1 * 2**-819:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0CC0000000000000;

    #10 $display("\n1 * 2**-820:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0CB0000000000000;

    #10 $display("\n1 * 2**-821:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0CA0000000000000;

    #10 $display("\n1 * 2**-822:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0C90000000000000;

    #10 $display("\n1 * 2**-823:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0C80000000000000;

    #10 $display("\n1 * 2**-824:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0C70000000000000;

    #10 $display("\n1 * 2**-825:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0C60000000000000;

    #10 $display("\n1 * 2**-826:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0C50000000000000;

    #10 $display("\n1 * 2**-827:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0C40000000000000;

    #10 $display("\n1 * 2**-828:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0C30000000000000;

    #10 $display("\n1 * 2**-829:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0C20000000000000;

    #10 $display("\n1 * 2**-830:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0C10000000000000;

    #10 $display("\n1 * 2**-831:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0C00000000000000;

    #10 $display("\n1 * 2**-832:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0BF0000000000000;

    #10 $display("\n1 * 2**-833:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0BE0000000000000;

    #10 $display("\n1 * 2**-834:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0BD0000000000000;

    #10 $display("\n1 * 2**-835:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0BC0000000000000;

    #10 $display("\n1 * 2**-836:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0BB0000000000000;

    #10 $display("\n1 * 2**-837:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0BA0000000000000;

    #10 $display("\n1 * 2**-838:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0B90000000000000;

    #10 $display("\n1 * 2**-839:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0B80000000000000;

    #10 $display("\n1 * 2**-840:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0B70000000000000;

    #10 $display("\n1 * 2**-841:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0B60000000000000;

    #10 $display("\n1 * 2**-842:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0B50000000000000;

    #10 $display("\n1 * 2**-843:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0B40000000000000;

    #10 $display("\n1 * 2**-844:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0B30000000000000;

    #10 $display("\n1 * 2**-845:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0B20000000000000;

    #10 $display("\n1 * 2**-846:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0B10000000000000;

    #10 $display("\n1 * 2**-847:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0B00000000000000;

    #10 $display("\n1 * 2**-848:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0AF0000000000000;

    #10 $display("\n1 * 2**-849:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0AE0000000000000;

    #10 $display("\n1 * 2**-850:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0AD0000000000000;

    #10 $display("\n1 * 2**-851:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0AC0000000000000;

    #10 $display("\n1 * 2**-852:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0AB0000000000000;

    #10 $display("\n1 * 2**-853:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0AA0000000000000;

    #10 $display("\n1 * 2**-854:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0A90000000000000;

    #10 $display("\n1 * 2**-855:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0A80000000000000;

    #10 $display("\n1 * 2**-856:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0A70000000000000;

    #10 $display("\n1 * 2**-857:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0A60000000000000;

    #10 $display("\n1 * 2**-858:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0A50000000000000;

    #10 $display("\n1 * 2**-859:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0A40000000000000;

    #10 $display("\n1 * 2**-860:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0A30000000000000;

    #10 $display("\n1 * 2**-861:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0A20000000000000;

    #10 $display("\n1 * 2**-862:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0A10000000000000;

    #10 $display("\n1 * 2**-863:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0A00000000000000;

    #10 $display("\n1 * 2**-864:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h09F0000000000000;

    #10 $display("\n1 * 2**-865:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h09E0000000000000;

    #10 $display("\n1 * 2**-866:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h09D0000000000000;

    #10 $display("\n1 * 2**-867:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h09C0000000000000;

    #10 $display("\n1 * 2**-868:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h09B0000000000000;

    #10 $display("\n1 * 2**-869:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h09A0000000000000;

    #10 $display("\n1 * 2**-870:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0990000000000000;

    #10 $display("\n1 * 2**-871:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0980000000000000;

    #10 $display("\n1 * 2**-872:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0970000000000000;

    #10 $display("\n1 * 2**-873:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0960000000000000;

    #10 $display("\n1 * 2**-874:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0950000000000000;

    #10 $display("\n1 * 2**-875:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0940000000000000;

    #10 $display("\n1 * 2**-876:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0930000000000000;

    #10 $display("\n1 * 2**-877:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0920000000000000;

    #10 $display("\n1 * 2**-878:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0910000000000000;

    #10 $display("\n1 * 2**-879:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0900000000000000;

    #10 $display("\n1 * 2**-880:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h08F0000000000000;

    #10 $display("\n1 * 2**-881:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h08E0000000000000;

    #10 $display("\n1 * 2**-882:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h08D0000000000000;

    #10 $display("\n1 * 2**-883:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h08C0000000000000;

    #10 $display("\n1 * 2**-884:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h08B0000000000000;

    #10 $display("\n1 * 2**-885:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h08A0000000000000;

    #10 $display("\n1 * 2**-886:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0890000000000000;

    #10 $display("\n1 * 2**-887:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0880000000000000;

    #10 $display("\n1 * 2**-888:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0870000000000000;

    #10 $display("\n1 * 2**-889:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0860000000000000;

    #10 $display("\n1 * 2**-890:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0850000000000000;

    #10 $display("\n1 * 2**-891:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0840000000000000;

    #10 $display("\n1 * 2**-892:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0830000000000000;

    #10 $display("\n1 * 2**-893:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0820000000000000;

    #10 $display("\n1 * 2**-894:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0810000000000000;

    #10 $display("\n1 * 2**-895:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0800000000000000;

    #10 $display("\n1 * 2**-896:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h07F0000000000000;

    #10 $display("\n1 * 2**-897:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h07E0000000000000;

    #10 $display("\n1 * 2**-898:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h07D0000000000000;

    #10 $display("\n1 * 2**-899:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h07C0000000000000;

    #10 $display("\n1 * 2**-900:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h07B0000000000000;

    #10 $display("\n1 * 2**-901:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h07A0000000000000;

    #10 $display("\n1 * 2**-902:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0790000000000000;

    #10 $display("\n1 * 2**-903:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0780000000000000;

    #10 $display("\n1 * 2**-904:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0770000000000000;

    #10 $display("\n1 * 2**-905:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0760000000000000;

    #10 $display("\n1 * 2**-906:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0750000000000000;

    #10 $display("\n1 * 2**-907:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0740000000000000;

    #10 $display("\n1 * 2**-908:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0730000000000000;

    #10 $display("\n1 * 2**-909:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0720000000000000;

    #10 $display("\n1 * 2**-910:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0710000000000000;

    #10 $display("\n1 * 2**-911:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0700000000000000;

    #10 $display("\n1 * 2**-912:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h06F0000000000000;

    #10 $display("\n1 * 2**-913:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h06E0000000000000;

    #10 $display("\n1 * 2**-914:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h06D0000000000000;

    #10 $display("\n1 * 2**-915:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h06C0000000000000;

    #10 $display("\n1 * 2**-916:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h06B0000000000000;

    #10 $display("\n1 * 2**-917:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h06A0000000000000;

    #10 $display("\n1 * 2**-918:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0690000000000000;

    #10 $display("\n1 * 2**-919:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0680000000000000;

    #10 $display("\n1 * 2**-920:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0670000000000000;

    #10 $display("\n1 * 2**-921:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0660000000000000;

    #10 $display("\n1 * 2**-922:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0650000000000000;

    #10 $display("\n1 * 2**-923:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0640000000000000;

    #10 $display("\n1 * 2**-924:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0630000000000000;

    #10 $display("\n1 * 2**-925:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0620000000000000;

    #10 $display("\n1 * 2**-926:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0610000000000000;

    #10 $display("\n1 * 2**-927:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0600000000000000;

    #10 $display("\n1 * 2**-928:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h05F0000000000000;

    #10 $display("\n1 * 2**-929:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h05E0000000000000;

    #10 $display("\n1 * 2**-930:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h05D0000000000000;

    #10 $display("\n1 * 2**-931:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h05C0000000000000;

    #10 $display("\n1 * 2**-932:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h05B0000000000000;

    #10 $display("\n1 * 2**-933:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h05A0000000000000;

    #10 $display("\n1 * 2**-934:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0590000000000000;

    #10 $display("\n1 * 2**-935:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0580000000000000;

    #10 $display("\n1 * 2**-936:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0570000000000000;

    #10 $display("\n1 * 2**-937:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0560000000000000;

    #10 $display("\n1 * 2**-938:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0550000000000000;

    #10 $display("\n1 * 2**-939:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0540000000000000;

    #10 $display("\n1 * 2**-940:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0530000000000000;

    #10 $display("\n1 * 2**-941:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0520000000000000;

    #10 $display("\n1 * 2**-942:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0510000000000000;

    #10 $display("\n1 * 2**-943:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0500000000000000;

    #10 $display("\n1 * 2**-944:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h04F0000000000000;

    #10 $display("\n1 * 2**-945:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h04E0000000000000;

    #10 $display("\n1 * 2**-946:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h04D0000000000000;

    #10 $display("\n1 * 2**-947:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h04C0000000000000;

    #10 $display("\n1 * 2**-948:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h04B0000000000000;

    #10 $display("\n1 * 2**-949:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h04A0000000000000;

    #10 $display("\n1 * 2**-950:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0490000000000000;

    #10 $display("\n1 * 2**-951:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0480000000000000;

    #10 $display("\n1 * 2**-952:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0470000000000000;

    #10 $display("\n1 * 2**-953:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0460000000000000;

    #10 $display("\n1 * 2**-954:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0450000000000000;

    #10 $display("\n1 * 2**-955:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0440000000000000;

    #10 $display("\n1 * 2**-956:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0430000000000000;

    #10 $display("\n1 * 2**-957:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0420000000000000;

    #10 $display("\n1 * 2**-958:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0410000000000000;

    #10 $display("\n1 * 2**-959:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0400000000000000;

    #10 $display("\n1 * 2**-960:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h03F0000000000000;

    #10 $display("\n1 * 2**-961:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h03E0000000000000;

    #10 $display("\n1 * 2**-962:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h03D0000000000000;

    #10 $display("\n1 * 2**-963:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h03C0000000000000;

    #10 $display("\n1 * 2**-964:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h03B0000000000000;

    #10 $display("\n1 * 2**-965:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h03A0000000000000;

    #10 $display("\n1 * 2**-966:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0390000000000000;

    #10 $display("\n1 * 2**-967:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0380000000000000;

    #10 $display("\n1 * 2**-968:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0370000000000000;

    #10 $display("\n1 * 2**-969:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0360000000000000;

    #10 $display("\n1 * 2**-970:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0350000000000000;

    #10 $display("\n1 * 2**-971:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0340000000000000;

    #10 $display("\n1 * 2**-972:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0330000000000000;

    #10 $display("\n1 * 2**-973:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0320000000000000;

    #10 $display("\n1 * 2**-974:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0310000000000000;

    #10 $display("\n1 * 2**-975:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0300000000000000;

    #10 $display("\n1 * 2**-976:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h02F0000000000000;

    #10 $display("\n1 * 2**-977:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h02E0000000000000;

    #10 $display("\n1 * 2**-978:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h02D0000000000000;

    #10 $display("\n1 * 2**-979:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h02C0000000000000;

    #10 $display("\n1 * 2**-980:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h02B0000000000000;

    #10 $display("\n1 * 2**-981:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h02A0000000000000;

    #10 $display("\n1 * 2**-982:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0290000000000000;

    #10 $display("\n1 * 2**-983:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0280000000000000;

    #10 $display("\n1 * 2**-984:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0270000000000000;

    #10 $display("\n1 * 2**-985:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0260000000000000;

    #10 $display("\n1 * 2**-986:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0250000000000000;

    #10 $display("\n1 * 2**-987:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0240000000000000;

    #10 $display("\n1 * 2**-988:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0230000000000000;

    #10 $display("\n1 * 2**-989:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0220000000000000;

    #10 $display("\n1 * 2**-990:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0210000000000000;

    #10 $display("\n1 * 2**-991:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0200000000000000;

    #10 $display("\n1 * 2**-992:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h01F0000000000000;

    #10 $display("\n1 * 2**-993:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h01E0000000000000;

    #10 $display("\n1 * 2**-994:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h01D0000000000000;

    #10 $display("\n1 * 2**-995:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h01C0000000000000;

    #10 $display("\n1 * 2**-996:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h01B0000000000000;

    #10 $display("\n1 * 2**-997:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h01A0000000000000;

    #10 $display("\n1 * 2**-998:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0190000000000000;

    #10 $display("\n1 * 2**-999:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0180000000000000;

    #10 $display("\n1 * 2**-1000:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0170000000000000;

    #10 $display("\n1 * 2**-1001:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0160000000000000;

    #10 $display("\n1 * 2**-1002:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0150000000000000;

    #10 $display("\n1 * 2**-1003:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0140000000000000;

    #10 $display("\n1 * 2**-1004:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0130000000000000;

    #10 $display("\n1 * 2**-1005:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0120000000000000;

    #10 $display("\n1 * 2**-1006:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0110000000000000;

    #10 $display("\n1 * 2**-1007:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0100000000000000;

    #10 $display("\n1 * 2**-1008:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h00F0000000000000;

    #10 $display("\n1 * 2**-1009:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h00E0000000000000;

    #10 $display("\n1 * 2**-1010:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h00D0000000000000;

    #10 $display("\n1 * 2**-1011:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h00C0000000000000;

    #10 $display("\n1 * 2**-1012:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h00B0000000000000;

    #10 $display("\n1 * 2**-1013:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h00A0000000000000;

    #10 $display("\n1 * 2**-1014:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0090000000000000;

    #10 $display("\n1 * 2**-1015:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0080000000000000;

    #10 $display("\n1 * 2**-1016:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0070000000000000;

    #10 $display("\n1 * 2**-1017:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0060000000000000;

    #10 $display("\n1 * 2**-1018:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0050000000000000;

    #10 $display("\n1 * 2**-1019:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0040000000000000;

    #10 $display("\n1 * 2**-1020:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0030000000000000;

    #10 $display("\n1 * 2**-1021:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0020000000000000;

    #10 $display("\n1 * 2**-1022:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0010000000000000;

    #10 $display("\n1 * 2**-1023:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0008000000000000;

    #10 $display("\n1 * 2**-1024:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0004000000000000;

    #10 $display("\n1 * 2**-1025:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0002000000000000;

    #10 $display("\n1 * 2**-1026:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0001000000000000;

    #10 $display("\n1 * 2**-1027:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000800000000000;

    #10 $display("\n1 * 2**-1028:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000400000000000;

    #10 $display("\n1 * 2**-1029:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000200000000000;

    #10 $display("\n1 * 2**-1030:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000100000000000;

    #10 $display("\n1 * 2**-1031:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000080000000000;

    #10 $display("\n1 * 2**-1032:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000040000000000;

    #10 $display("\n1 * 2**-1033:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000020000000000;

    #10 $display("\n1 * 2**-1034:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000010000000000;

    #10 $display("\n1 * 2**-1035:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000008000000000;

    #10 $display("\n1 * 2**-1036:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000004000000000;

    #10 $display("\n1 * 2**-1037:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000002000000000;

    #10 $display("\n1 * 2**-1038:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000001000000000;

    #10 $display("\n1 * 2**-1039:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000800000000;

    #10 $display("\n1 * 2**-1040:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000400000000;

    #10 $display("\n1 * 2**-1041:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000200000000;

    #10 $display("\n1 * 2**-1042:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000100000000;

    #10 $display("\n1 * 2**-1043:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000080000000;

    #10 $display("\n1 * 2**-1044:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000040000000;

    #10 $display("\n1 * 2**-1045:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000020000000;

    #10 $display("\n1 * 2**-1046:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000010000000;

    #10 $display("\n1 * 2**-1047:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000008000000;

    #10 $display("\n1 * 2**-1048:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000004000000;

    #10 $display("\n1 * 2**-1049:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000002000000;

    #10 $display("\n1 * 2**-1050:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000001000000;

    #10 $display("\n1 * 2**-1051:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000800000;

    #10 $display("\n1 * 2**-1052:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000400000;

    #10 $display("\n1 * 2**-1053:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000200000;

    #10 $display("\n1 * 2**-1054:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000100000;

    #10 $display("\n1 * 2**-1055:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000080000;

    #10 $display("\n1 * 2**-1056:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000040000;

    #10 $display("\n1 * 2**-1057:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000020000;

    #10 $display("\n1 * 2**-1058:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000010000;

    #10 $display("\n1 * 2**-1059:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000008000;

    #10 $display("\n1 * 2**-1060:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000004000;

    #10 $display("\n1 * 2**-1061:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000002000;

    #10 $display("\n1 * 2**-1062:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000001000;

    #10 $display("\n1 * 2**-1063:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000000800;

    #10 $display("\n1 * 2**-1064:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000000400;

    #10 $display("\n1 * 2**-1065:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000000200;

    #10 $display("\n1 * 2**-1066:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000000100;

    #10 $display("\n1 * 2**-1067:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000000080;

    #10 $display("\n1 * 2**-1068:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000000040;

    #10 $display("\n1 * 2**-1069:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000000020;

    #10 $display("\n1 * 2**-1070:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000000010;

    #10 $display("\n1 * 2**-1071:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000000008;

    #10 $display("\n1 * 2**-1072:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000000004;

    #10 $display("\n1 * 2**-1073:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000000002;

    #10 $display("\n1 * 2**-1074:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0000000000000001;

    #10 $display("\n2**1023 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7FE0000000000000;

    #10 $display("\n2**1022 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7FD0000000000000;

    #10 $display("\n2**1021 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7FC0000000000000;

    #10 $display("\n2**1020 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7FB0000000000000;

    #10 $display("\n2**1019 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7FA0000000000000;

    #10 $display("\n2**1018 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7F90000000000000;

    #10 $display("\n2**1017 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7F80000000000000;

    #10 $display("\n2**1016 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7F70000000000000;

    #10 $display("\n2**1015 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7F60000000000000;

    #10 $display("\n2**1014 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7F50000000000000;

    #10 $display("\n2**1013 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7F40000000000000;

    #10 $display("\n2**1012 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7F30000000000000;

    #10 $display("\n2**1011 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7F20000000000000;

    #10 $display("\n2**1010 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7F10000000000000;

    #10 $display("\n2**1009 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7F00000000000000;

    #10 $display("\n2**1008 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7EF0000000000000;

    #10 $display("\n2**1007 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7EE0000000000000;

    #10 $display("\n2**1006 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7ED0000000000000;

    #10 $display("\n2**1005 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7EC0000000000000;

    #10 $display("\n2**1004 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7EB0000000000000;

    #10 $display("\n2**1003 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7EA0000000000000;

    #10 $display("\n2**1002 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7E90000000000000;

    #10 $display("\n2**1001 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7E80000000000000;

    #10 $display("\n2**1000 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7E70000000000000;

    #10 $display("\n2**999 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7E60000000000000;

    #10 $display("\n2**998 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7E50000000000000;

    #10 $display("\n2**997 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7E40000000000000;

    #10 $display("\n2**996 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7E30000000000000;

    #10 $display("\n2**995 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7E20000000000000;

    #10 $display("\n2**994 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7E10000000000000;

    #10 $display("\n2**993 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7E00000000000000;

    #10 $display("\n2**992 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7DF0000000000000;

    #10 $display("\n2**991 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7DE0000000000000;

    #10 $display("\n2**990 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7DD0000000000000;

    #10 $display("\n2**989 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7DC0000000000000;

    #10 $display("\n2**988 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7DB0000000000000;

    #10 $display("\n2**987 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7DA0000000000000;

    #10 $display("\n2**986 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7D90000000000000;

    #10 $display("\n2**985 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7D80000000000000;

    #10 $display("\n2**984 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7D70000000000000;

    #10 $display("\n2**983 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7D60000000000000;

    #10 $display("\n2**982 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7D50000000000000;

    #10 $display("\n2**981 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7D40000000000000;

    #10 $display("\n2**980 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7D30000000000000;

    #10 $display("\n2**979 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7D20000000000000;

    #10 $display("\n2**978 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7D10000000000000;

    #10 $display("\n2**977 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7D00000000000000;

    #10 $display("\n2**976 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7CF0000000000000;

    #10 $display("\n2**975 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7CE0000000000000;

    #10 $display("\n2**974 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7CD0000000000000;

    #10 $display("\n2**973 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7CC0000000000000;

    #10 $display("\n2**972 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7CB0000000000000;

    #10 $display("\n2**971 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7CA0000000000000;

    #10 $display("\n2**970 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7C90000000000000;

    #10 $display("\n2**969 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7C80000000000000;

    #10 $display("\n2**968 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7C70000000000000;

    #10 $display("\n2**967 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7C60000000000000;

    #10 $display("\n2**966 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7C50000000000000;

    #10 $display("\n2**965 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7C40000000000000;

    #10 $display("\n2**964 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7C30000000000000;

    #10 $display("\n2**963 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7C20000000000000;

    #10 $display("\n2**962 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7C10000000000000;

    #10 $display("\n2**961 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7C00000000000000;

    #10 $display("\n2**960 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7BF0000000000000;

    #10 $display("\n2**959 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7BE0000000000000;

    #10 $display("\n2**958 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7BD0000000000000;

    #10 $display("\n2**957 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7BC0000000000000;

    #10 $display("\n2**956 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7BB0000000000000;

    #10 $display("\n2**955 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7BA0000000000000;

    #10 $display("\n2**954 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7B90000000000000;

    #10 $display("\n2**953 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7B80000000000000;

    #10 $display("\n2**952 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7B70000000000000;

    #10 $display("\n2**951 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7B60000000000000;

    #10 $display("\n2**950 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7B50000000000000;

    #10 $display("\n2**949 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7B40000000000000;

    #10 $display("\n2**948 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7B30000000000000;

    #10 $display("\n2**947 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7B20000000000000;

    #10 $display("\n2**946 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7B10000000000000;

    #10 $display("\n2**945 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7B00000000000000;

    #10 $display("\n2**944 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7AF0000000000000;

    #10 $display("\n2**943 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7AE0000000000000;

    #10 $display("\n2**942 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7AD0000000000000;

    #10 $display("\n2**941 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7AC0000000000000;

    #10 $display("\n2**940 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7AB0000000000000;

    #10 $display("\n2**939 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7AA0000000000000;

    #10 $display("\n2**938 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7A90000000000000;

    #10 $display("\n2**937 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7A80000000000000;

    #10 $display("\n2**936 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7A70000000000000;

    #10 $display("\n2**935 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7A60000000000000;

    #10 $display("\n2**934 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7A50000000000000;

    #10 $display("\n2**933 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7A40000000000000;

    #10 $display("\n2**932 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7A30000000000000;

    #10 $display("\n2**931 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7A20000000000000;

    #10 $display("\n2**930 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7A10000000000000;

    #10 $display("\n2**929 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7A00000000000000;

    #10 $display("\n2**928 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h79F0000000000000;

    #10 $display("\n2**927 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h79E0000000000000;

    #10 $display("\n2**926 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h79D0000000000000;

    #10 $display("\n2**925 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h79C0000000000000;

    #10 $display("\n2**924 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h79B0000000000000;

    #10 $display("\n2**923 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h79A0000000000000;

    #10 $display("\n2**922 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7990000000000000;

    #10 $display("\n2**921 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7980000000000000;

    #10 $display("\n2**920 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7970000000000000;

    #10 $display("\n2**919 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7960000000000000;

    #10 $display("\n2**918 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7950000000000000;

    #10 $display("\n2**917 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7940000000000000;

    #10 $display("\n2**916 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7930000000000000;

    #10 $display("\n2**915 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7920000000000000;

    #10 $display("\n2**914 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7910000000000000;

    #10 $display("\n2**913 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7900000000000000;

    #10 $display("\n2**912 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h78F0000000000000;

    #10 $display("\n2**911 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h78E0000000000000;

    #10 $display("\n2**910 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h78D0000000000000;

    #10 $display("\n2**909 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h78C0000000000000;

    #10 $display("\n2**908 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h78B0000000000000;

    #10 $display("\n2**907 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h78A0000000000000;

    #10 $display("\n2**906 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7890000000000000;

    #10 $display("\n2**905 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7880000000000000;

    #10 $display("\n2**904 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7870000000000000;

    #10 $display("\n2**903 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7860000000000000;

    #10 $display("\n2**902 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7850000000000000;

    #10 $display("\n2**901 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7840000000000000;

    #10 $display("\n2**900 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7830000000000000;

    #10 $display("\n2**899 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7820000000000000;

    #10 $display("\n2**898 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7810000000000000;

    #10 $display("\n2**897 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7800000000000000;

    #10 $display("\n2**896 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h77F0000000000000;

    #10 $display("\n2**895 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h77E0000000000000;

    #10 $display("\n2**894 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h77D0000000000000;

    #10 $display("\n2**893 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h77C0000000000000;

    #10 $display("\n2**892 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h77B0000000000000;

    #10 $display("\n2**891 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h77A0000000000000;

    #10 $display("\n2**890 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7790000000000000;

    #10 $display("\n2**889 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7780000000000000;

    #10 $display("\n2**888 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7770000000000000;

    #10 $display("\n2**887 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7760000000000000;

    #10 $display("\n2**886 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7750000000000000;

    #10 $display("\n2**885 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7740000000000000;

    #10 $display("\n2**884 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7730000000000000;

    #10 $display("\n2**883 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7720000000000000;

    #10 $display("\n2**882 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7710000000000000;

    #10 $display("\n2**881 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7700000000000000;

    #10 $display("\n2**880 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h76F0000000000000;

    #10 $display("\n2**879 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h76E0000000000000;

    #10 $display("\n2**878 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h76D0000000000000;

    #10 $display("\n2**877 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h76C0000000000000;

    #10 $display("\n2**876 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h76B0000000000000;

    #10 $display("\n2**875 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h76A0000000000000;

    #10 $display("\n2**874 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7690000000000000;

    #10 $display("\n2**873 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7680000000000000;

    #10 $display("\n2**872 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7670000000000000;

    #10 $display("\n2**871 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7660000000000000;

    #10 $display("\n2**870 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7650000000000000;

    #10 $display("\n2**869 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7640000000000000;

    #10 $display("\n2**868 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7630000000000000;

    #10 $display("\n2**867 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7620000000000000;

    #10 $display("\n2**866 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7610000000000000;

    #10 $display("\n2**865 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7600000000000000;

    #10 $display("\n2**864 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h75F0000000000000;

    #10 $display("\n2**863 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h75E0000000000000;

    #10 $display("\n2**862 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h75D0000000000000;

    #10 $display("\n2**861 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h75C0000000000000;

    #10 $display("\n2**860 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h75B0000000000000;

    #10 $display("\n2**859 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h75A0000000000000;

    #10 $display("\n2**858 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7590000000000000;

    #10 $display("\n2**857 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7580000000000000;

    #10 $display("\n2**856 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7570000000000000;

    #10 $display("\n2**855 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7560000000000000;

    #10 $display("\n2**854 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7550000000000000;

    #10 $display("\n2**853 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7540000000000000;

    #10 $display("\n2**852 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7530000000000000;

    #10 $display("\n2**851 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7520000000000000;

    #10 $display("\n2**850 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7510000000000000;

    #10 $display("\n2**849 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7500000000000000;

    #10 $display("\n2**848 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h74F0000000000000;

    #10 $display("\n2**847 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h74E0000000000000;

    #10 $display("\n2**846 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h74D0000000000000;

    #10 $display("\n2**845 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h74C0000000000000;

    #10 $display("\n2**844 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h74B0000000000000;

    #10 $display("\n2**843 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h74A0000000000000;

    #10 $display("\n2**842 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7490000000000000;

    #10 $display("\n2**841 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7480000000000000;

    #10 $display("\n2**840 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7470000000000000;

    #10 $display("\n2**839 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7460000000000000;

    #10 $display("\n2**838 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7450000000000000;

    #10 $display("\n2**837 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7440000000000000;

    #10 $display("\n2**836 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7430000000000000;

    #10 $display("\n2**835 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7420000000000000;

    #10 $display("\n2**834 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7410000000000000;

    #10 $display("\n2**833 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7400000000000000;

    #10 $display("\n2**832 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h73F0000000000000;

    #10 $display("\n2**831 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h73E0000000000000;

    #10 $display("\n2**830 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h73D0000000000000;

    #10 $display("\n2**829 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h73C0000000000000;

    #10 $display("\n2**828 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h73B0000000000000;

    #10 $display("\n2**827 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h73A0000000000000;

    #10 $display("\n2**826 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7390000000000000;

    #10 $display("\n2**825 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7380000000000000;

    #10 $display("\n2**824 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7370000000000000;

    #10 $display("\n2**823 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7360000000000000;

    #10 $display("\n2**822 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7350000000000000;

    #10 $display("\n2**821 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7340000000000000;

    #10 $display("\n2**820 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7330000000000000;

    #10 $display("\n2**819 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7320000000000000;

    #10 $display("\n2**818 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7310000000000000;

    #10 $display("\n2**817 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7300000000000000;

    #10 $display("\n2**816 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h72F0000000000000;

    #10 $display("\n2**815 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h72E0000000000000;

    #10 $display("\n2**814 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h72D0000000000000;

    #10 $display("\n2**813 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h72C0000000000000;

    #10 $display("\n2**812 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h72B0000000000000;

    #10 $display("\n2**811 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h72A0000000000000;

    #10 $display("\n2**810 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7290000000000000;

    #10 $display("\n2**809 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7280000000000000;

    #10 $display("\n2**808 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7270000000000000;

    #10 $display("\n2**807 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7260000000000000;

    #10 $display("\n2**806 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7250000000000000;

    #10 $display("\n2**805 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7240000000000000;

    #10 $display("\n2**804 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7230000000000000;

    #10 $display("\n2**803 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7220000000000000;

    #10 $display("\n2**802 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7210000000000000;

    #10 $display("\n2**801 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7200000000000000;

    #10 $display("\n2**800 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h71F0000000000000;

    #10 $display("\n2**799 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h71E0000000000000;

    #10 $display("\n2**798 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h71D0000000000000;

    #10 $display("\n2**797 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h71C0000000000000;

    #10 $display("\n2**796 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h71B0000000000000;

    #10 $display("\n2**795 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h71A0000000000000;

    #10 $display("\n2**794 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7190000000000000;

    #10 $display("\n2**793 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7180000000000000;

    #10 $display("\n2**792 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7170000000000000;

    #10 $display("\n2**791 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7160000000000000;

    #10 $display("\n2**790 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7150000000000000;

    #10 $display("\n2**789 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7140000000000000;

    #10 $display("\n2**788 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7130000000000000;

    #10 $display("\n2**787 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7120000000000000;

    #10 $display("\n2**786 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7110000000000000;

    #10 $display("\n2**785 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7100000000000000;

    #10 $display("\n2**784 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h70F0000000000000;

    #10 $display("\n2**783 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h70E0000000000000;

    #10 $display("\n2**782 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h70D0000000000000;

    #10 $display("\n2**781 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h70C0000000000000;

    #10 $display("\n2**780 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h70B0000000000000;

    #10 $display("\n2**779 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h70A0000000000000;

    #10 $display("\n2**778 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7090000000000000;

    #10 $display("\n2**777 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7080000000000000;

    #10 $display("\n2**776 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7070000000000000;

    #10 $display("\n2**775 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7060000000000000;

    #10 $display("\n2**774 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7050000000000000;

    #10 $display("\n2**773 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7040000000000000;

    #10 $display("\n2**772 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7030000000000000;

    #10 $display("\n2**771 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7020000000000000;

    #10 $display("\n2**770 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7010000000000000;

    #10 $display("\n2**769 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h7000000000000000;

    #10 $display("\n2**768 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6FF0000000000000;

    #10 $display("\n2**767 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6FE0000000000000;

    #10 $display("\n2**766 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6FD0000000000000;

    #10 $display("\n2**765 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6FC0000000000000;

    #10 $display("\n2**764 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6FB0000000000000;

    #10 $display("\n2**763 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6FA0000000000000;

    #10 $display("\n2**762 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6F90000000000000;

    #10 $display("\n2**761 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6F80000000000000;

    #10 $display("\n2**760 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6F70000000000000;

    #10 $display("\n2**759 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6F60000000000000;

    #10 $display("\n2**758 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6F50000000000000;

    #10 $display("\n2**757 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6F40000000000000;

    #10 $display("\n2**756 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6F30000000000000;

    #10 $display("\n2**755 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6F20000000000000;

    #10 $display("\n2**754 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6F10000000000000;

    #10 $display("\n2**753 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6F00000000000000;

    #10 $display("\n2**752 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6EF0000000000000;

    #10 $display("\n2**751 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6EE0000000000000;

    #10 $display("\n2**750 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6ED0000000000000;

    #10 $display("\n2**749 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6EC0000000000000;

    #10 $display("\n2**748 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6EB0000000000000;

    #10 $display("\n2**747 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6EA0000000000000;

    #10 $display("\n2**746 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6E90000000000000;

    #10 $display("\n2**745 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6E80000000000000;

    #10 $display("\n2**744 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6E70000000000000;

    #10 $display("\n2**743 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6E60000000000000;

    #10 $display("\n2**742 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6E50000000000000;

    #10 $display("\n2**741 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6E40000000000000;

    #10 $display("\n2**740 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6E30000000000000;

    #10 $display("\n2**739 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6E20000000000000;

    #10 $display("\n2**738 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6E10000000000000;

    #10 $display("\n2**737 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6E00000000000000;

    #10 $display("\n2**736 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6DF0000000000000;

    #10 $display("\n2**735 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6DE0000000000000;

    #10 $display("\n2**734 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6DD0000000000000;

    #10 $display("\n2**733 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6DC0000000000000;

    #10 $display("\n2**732 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6DB0000000000000;

    #10 $display("\n2**731 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6DA0000000000000;

    #10 $display("\n2**730 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6D90000000000000;

    #10 $display("\n2**729 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6D80000000000000;

    #10 $display("\n2**728 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6D70000000000000;

    #10 $display("\n2**727 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6D60000000000000;

    #10 $display("\n2**726 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6D50000000000000;

    #10 $display("\n2**725 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6D40000000000000;

    #10 $display("\n2**724 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6D30000000000000;

    #10 $display("\n2**723 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6D20000000000000;

    #10 $display("\n2**722 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6D10000000000000;

    #10 $display("\n2**721 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6D00000000000000;

    #10 $display("\n2**720 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6CF0000000000000;

    #10 $display("\n2**719 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6CE0000000000000;

    #10 $display("\n2**718 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6CD0000000000000;

    #10 $display("\n2**717 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6CC0000000000000;

    #10 $display("\n2**716 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6CB0000000000000;

    #10 $display("\n2**715 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6CA0000000000000;

    #10 $display("\n2**714 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6C90000000000000;

    #10 $display("\n2**713 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6C80000000000000;

    #10 $display("\n2**712 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6C70000000000000;

    #10 $display("\n2**711 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6C60000000000000;

    #10 $display("\n2**710 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6C50000000000000;

    #10 $display("\n2**709 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6C40000000000000;

    #10 $display("\n2**708 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6C30000000000000;

    #10 $display("\n2**707 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6C20000000000000;

    #10 $display("\n2**706 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6C10000000000000;

    #10 $display("\n2**705 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6C00000000000000;

    #10 $display("\n2**704 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6BF0000000000000;

    #10 $display("\n2**703 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6BE0000000000000;

    #10 $display("\n2**702 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6BD0000000000000;

    #10 $display("\n2**701 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6BC0000000000000;

    #10 $display("\n2**700 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6BB0000000000000;

    #10 $display("\n2**699 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6BA0000000000000;

    #10 $display("\n2**698 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6B90000000000000;

    #10 $display("\n2**697 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6B80000000000000;

    #10 $display("\n2**696 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6B70000000000000;

    #10 $display("\n2**695 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6B60000000000000;

    #10 $display("\n2**694 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6B50000000000000;

    #10 $display("\n2**693 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6B40000000000000;

    #10 $display("\n2**692 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6B30000000000000;

    #10 $display("\n2**691 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6B20000000000000;

    #10 $display("\n2**690 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6B10000000000000;

    #10 $display("\n2**689 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6B00000000000000;

    #10 $display("\n2**688 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6AF0000000000000;

    #10 $display("\n2**687 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6AE0000000000000;

    #10 $display("\n2**686 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6AD0000000000000;

    #10 $display("\n2**685 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6AC0000000000000;

    #10 $display("\n2**684 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6AB0000000000000;

    #10 $display("\n2**683 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6AA0000000000000;

    #10 $display("\n2**682 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6A90000000000000;

    #10 $display("\n2**681 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6A80000000000000;

    #10 $display("\n2**680 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6A70000000000000;

    #10 $display("\n2**679 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6A60000000000000;

    #10 $display("\n2**678 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6A50000000000000;

    #10 $display("\n2**677 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6A40000000000000;

    #10 $display("\n2**676 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6A30000000000000;

    #10 $display("\n2**675 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6A20000000000000;

    #10 $display("\n2**674 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6A10000000000000;

    #10 $display("\n2**673 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6A00000000000000;

    #10 $display("\n2**672 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h69F0000000000000;

    #10 $display("\n2**671 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h69E0000000000000;

    #10 $display("\n2**670 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h69D0000000000000;

    #10 $display("\n2**669 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h69C0000000000000;

    #10 $display("\n2**668 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h69B0000000000000;

    #10 $display("\n2**667 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h69A0000000000000;

    #10 $display("\n2**666 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6990000000000000;

    #10 $display("\n2**665 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6980000000000000;

    #10 $display("\n2**664 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6970000000000000;

    #10 $display("\n2**663 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6960000000000000;

    #10 $display("\n2**662 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6950000000000000;

    #10 $display("\n2**661 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6940000000000000;

    #10 $display("\n2**660 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6930000000000000;

    #10 $display("\n2**659 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6920000000000000;

    #10 $display("\n2**658 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6910000000000000;

    #10 $display("\n2**657 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6900000000000000;

    #10 $display("\n2**656 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h68F0000000000000;

    #10 $display("\n2**655 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h68E0000000000000;

    #10 $display("\n2**654 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h68D0000000000000;

    #10 $display("\n2**653 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h68C0000000000000;

    #10 $display("\n2**652 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h68B0000000000000;

    #10 $display("\n2**651 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h68A0000000000000;

    #10 $display("\n2**650 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6890000000000000;

    #10 $display("\n2**649 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6880000000000000;

    #10 $display("\n2**648 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6870000000000000;

    #10 $display("\n2**647 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6860000000000000;

    #10 $display("\n2**646 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6850000000000000;

    #10 $display("\n2**645 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6840000000000000;

    #10 $display("\n2**644 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6830000000000000;

    #10 $display("\n2**643 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6820000000000000;

    #10 $display("\n2**642 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6810000000000000;

    #10 $display("\n2**641 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6800000000000000;

    #10 $display("\n2**640 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h67F0000000000000;

    #10 $display("\n2**639 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h67E0000000000000;

    #10 $display("\n2**638 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h67D0000000000000;

    #10 $display("\n2**637 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h67C0000000000000;

    #10 $display("\n2**636 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h67B0000000000000;

    #10 $display("\n2**635 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h67A0000000000000;

    #10 $display("\n2**634 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6790000000000000;

    #10 $display("\n2**633 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6780000000000000;

    #10 $display("\n2**632 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6770000000000000;

    #10 $display("\n2**631 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6760000000000000;

    #10 $display("\n2**630 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6750000000000000;

    #10 $display("\n2**629 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6740000000000000;

    #10 $display("\n2**628 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6730000000000000;

    #10 $display("\n2**627 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6720000000000000;

    #10 $display("\n2**626 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6710000000000000;

    #10 $display("\n2**625 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6700000000000000;

    #10 $display("\n2**624 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h66F0000000000000;

    #10 $display("\n2**623 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h66E0000000000000;

    #10 $display("\n2**622 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h66D0000000000000;

    #10 $display("\n2**621 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h66C0000000000000;

    #10 $display("\n2**620 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h66B0000000000000;

    #10 $display("\n2**619 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h66A0000000000000;

    #10 $display("\n2**618 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6690000000000000;

    #10 $display("\n2**617 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6680000000000000;

    #10 $display("\n2**616 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6670000000000000;

    #10 $display("\n2**615 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6660000000000000;

    #10 $display("\n2**614 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6650000000000000;

    #10 $display("\n2**613 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6640000000000000;

    #10 $display("\n2**612 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6630000000000000;

    #10 $display("\n2**611 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6620000000000000;

    #10 $display("\n2**610 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6610000000000000;

    #10 $display("\n2**609 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6600000000000000;

    #10 $display("\n2**608 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h65F0000000000000;

    #10 $display("\n2**607 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h65E0000000000000;

    #10 $display("\n2**606 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h65D0000000000000;

    #10 $display("\n2**605 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h65C0000000000000;

    #10 $display("\n2**604 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h65B0000000000000;

    #10 $display("\n2**603 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h65A0000000000000;

    #10 $display("\n2**602 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6590000000000000;

    #10 $display("\n2**601 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6580000000000000;

    #10 $display("\n2**600 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6570000000000000;

    #10 $display("\n2**599 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6560000000000000;

    #10 $display("\n2**598 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6550000000000000;

    #10 $display("\n2**597 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6540000000000000;

    #10 $display("\n2**596 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6530000000000000;

    #10 $display("\n2**595 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6520000000000000;

    #10 $display("\n2**594 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6510000000000000;

    #10 $display("\n2**593 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6500000000000000;

    #10 $display("\n2**592 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h64F0000000000000;

    #10 $display("\n2**591 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h64E0000000000000;

    #10 $display("\n2**590 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h64D0000000000000;

    #10 $display("\n2**589 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h64C0000000000000;

    #10 $display("\n2**588 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h64B0000000000000;

    #10 $display("\n2**587 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h64A0000000000000;

    #10 $display("\n2**586 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6490000000000000;

    #10 $display("\n2**585 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6480000000000000;

    #10 $display("\n2**584 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6470000000000000;

    #10 $display("\n2**583 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6460000000000000;

    #10 $display("\n2**582 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6450000000000000;

    #10 $display("\n2**581 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6440000000000000;

    #10 $display("\n2**580 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6430000000000000;

    #10 $display("\n2**579 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6420000000000000;

    #10 $display("\n2**578 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6410000000000000;

    #10 $display("\n2**577 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6400000000000000;

    #10 $display("\n2**576 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h63F0000000000000;

    #10 $display("\n2**575 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h63E0000000000000;

    #10 $display("\n2**574 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h63D0000000000000;

    #10 $display("\n2**573 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h63C0000000000000;

    #10 $display("\n2**572 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h63B0000000000000;

    #10 $display("\n2**571 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h63A0000000000000;

    #10 $display("\n2**570 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6390000000000000;

    #10 $display("\n2**569 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6380000000000000;

    #10 $display("\n2**568 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6370000000000000;

    #10 $display("\n2**567 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6360000000000000;

    #10 $display("\n2**566 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6350000000000000;

    #10 $display("\n2**565 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6340000000000000;

    #10 $display("\n2**564 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6330000000000000;

    #10 $display("\n2**563 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6320000000000000;

    #10 $display("\n2**562 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6310000000000000;

    #10 $display("\n2**561 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6300000000000000;

    #10 $display("\n2**560 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h62F0000000000000;

    #10 $display("\n2**559 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h62E0000000000000;

    #10 $display("\n2**558 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h62D0000000000000;

    #10 $display("\n2**557 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h62C0000000000000;

    #10 $display("\n2**556 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h62B0000000000000;

    #10 $display("\n2**555 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h62A0000000000000;

    #10 $display("\n2**554 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6290000000000000;

    #10 $display("\n2**553 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6280000000000000;

    #10 $display("\n2**552 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6270000000000000;

    #10 $display("\n2**551 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6260000000000000;

    #10 $display("\n2**550 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6250000000000000;

    #10 $display("\n2**549 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6240000000000000;

    #10 $display("\n2**548 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6230000000000000;

    #10 $display("\n2**547 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6220000000000000;

    #10 $display("\n2**546 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6210000000000000;

    #10 $display("\n2**545 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6200000000000000;

    #10 $display("\n2**544 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h61F0000000000000;

    #10 $display("\n2**543 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h61E0000000000000;

    #10 $display("\n2**542 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h61D0000000000000;

    #10 $display("\n2**541 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h61C0000000000000;

    #10 $display("\n2**540 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h61B0000000000000;

    #10 $display("\n2**539 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h61A0000000000000;

    #10 $display("\n2**538 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6190000000000000;

    #10 $display("\n2**537 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6180000000000000;

    #10 $display("\n2**536 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6170000000000000;

    #10 $display("\n2**535 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6160000000000000;

    #10 $display("\n2**534 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6150000000000000;

    #10 $display("\n2**533 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6140000000000000;

    #10 $display("\n2**532 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6130000000000000;

    #10 $display("\n2**531 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6120000000000000;

    #10 $display("\n2**530 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6110000000000000;

    #10 $display("\n2**529 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6100000000000000;

    #10 $display("\n2**528 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h60F0000000000000;

    #10 $display("\n2**527 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h60E0000000000000;

    #10 $display("\n2**526 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h60D0000000000000;

    #10 $display("\n2**525 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h60C0000000000000;

    #10 $display("\n2**524 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h60B0000000000000;

    #10 $display("\n2**523 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h60A0000000000000;

    #10 $display("\n2**522 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6090000000000000;

    #10 $display("\n2**521 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6080000000000000;

    #10 $display("\n2**520 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6070000000000000;

    #10 $display("\n2**519 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6060000000000000;

    #10 $display("\n2**518 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6050000000000000;

    #10 $display("\n2**517 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6040000000000000;

    #10 $display("\n2**516 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6030000000000000;

    #10 $display("\n2**515 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6020000000000000;

    #10 $display("\n2**514 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6010000000000000;

    #10 $display("\n2**513 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h6000000000000000;

    #10 $display("\n2**512 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5FF0000000000000;

    #10 $display("\n2**511 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5FE0000000000000;

    #10 $display("\n2**510 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5FD0000000000000;

    #10 $display("\n2**509 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5FC0000000000000;

    #10 $display("\n2**508 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5FB0000000000000;

    #10 $display("\n2**507 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5FA0000000000000;

    #10 $display("\n2**506 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5F90000000000000;

    #10 $display("\n2**505 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5F80000000000000;

    #10 $display("\n2**504 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5F70000000000000;

    #10 $display("\n2**503 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5F60000000000000;

    #10 $display("\n2**502 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5F50000000000000;

    #10 $display("\n2**501 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5F40000000000000;

    #10 $display("\n2**500 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5F30000000000000;

    #10 $display("\n2**499 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5F20000000000000;

    #10 $display("\n2**498 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5F10000000000000;

    #10 $display("\n2**497 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5F00000000000000;

    #10 $display("\n2**496 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5EF0000000000000;

    #10 $display("\n2**495 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5EE0000000000000;

    #10 $display("\n2**494 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5ED0000000000000;

    #10 $display("\n2**493 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5EC0000000000000;

    #10 $display("\n2**492 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5EB0000000000000;

    #10 $display("\n2**491 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5EA0000000000000;

    #10 $display("\n2**490 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5E90000000000000;

    #10 $display("\n2**489 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5E80000000000000;

    #10 $display("\n2**488 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5E70000000000000;

    #10 $display("\n2**487 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5E60000000000000;

    #10 $display("\n2**486 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5E50000000000000;

    #10 $display("\n2**485 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5E40000000000000;

    #10 $display("\n2**484 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5E30000000000000;

    #10 $display("\n2**483 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5E20000000000000;

    #10 $display("\n2**482 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5E10000000000000;

    #10 $display("\n2**481 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5E00000000000000;

    #10 $display("\n2**480 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5DF0000000000000;

    #10 $display("\n2**479 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5DE0000000000000;

    #10 $display("\n2**478 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5DD0000000000000;

    #10 $display("\n2**477 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5DC0000000000000;

    #10 $display("\n2**476 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5DB0000000000000;

    #10 $display("\n2**475 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5DA0000000000000;

    #10 $display("\n2**474 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5D90000000000000;

    #10 $display("\n2**473 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5D80000000000000;

    #10 $display("\n2**472 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5D70000000000000;

    #10 $display("\n2**471 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5D60000000000000;

    #10 $display("\n2**470 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5D50000000000000;

    #10 $display("\n2**469 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5D40000000000000;

    #10 $display("\n2**468 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5D30000000000000;

    #10 $display("\n2**467 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5D20000000000000;

    #10 $display("\n2**466 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5D10000000000000;

    #10 $display("\n2**465 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5D00000000000000;

    #10 $display("\n2**464 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5CF0000000000000;

    #10 $display("\n2**463 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5CE0000000000000;

    #10 $display("\n2**462 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5CD0000000000000;

    #10 $display("\n2**461 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5CC0000000000000;

    #10 $display("\n2**460 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5CB0000000000000;

    #10 $display("\n2**459 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5CA0000000000000;

    #10 $display("\n2**458 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5C90000000000000;

    #10 $display("\n2**457 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5C80000000000000;

    #10 $display("\n2**456 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5C70000000000000;

    #10 $display("\n2**455 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5C60000000000000;

    #10 $display("\n2**454 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5C50000000000000;

    #10 $display("\n2**453 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5C40000000000000;

    #10 $display("\n2**452 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5C30000000000000;

    #10 $display("\n2**451 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5C20000000000000;

    #10 $display("\n2**450 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5C10000000000000;

    #10 $display("\n2**449 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5C00000000000000;

    #10 $display("\n2**448 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5BF0000000000000;

    #10 $display("\n2**447 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5BE0000000000000;

    #10 $display("\n2**446 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5BD0000000000000;

    #10 $display("\n2**445 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5BC0000000000000;

    #10 $display("\n2**444 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5BB0000000000000;

    #10 $display("\n2**443 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5BA0000000000000;

    #10 $display("\n2**442 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5B90000000000000;

    #10 $display("\n2**441 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5B80000000000000;

    #10 $display("\n2**440 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5B70000000000000;

    #10 $display("\n2**439 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5B60000000000000;

    #10 $display("\n2**438 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5B50000000000000;

    #10 $display("\n2**437 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5B40000000000000;

    #10 $display("\n2**436 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5B30000000000000;

    #10 $display("\n2**435 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5B20000000000000;

    #10 $display("\n2**434 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5B10000000000000;

    #10 $display("\n2**433 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5B00000000000000;

    #10 $display("\n2**432 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5AF0000000000000;

    #10 $display("\n2**431 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5AE0000000000000;

    #10 $display("\n2**430 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5AD0000000000000;

    #10 $display("\n2**429 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5AC0000000000000;

    #10 $display("\n2**428 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5AB0000000000000;

    #10 $display("\n2**427 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5AA0000000000000;

    #10 $display("\n2**426 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5A90000000000000;

    #10 $display("\n2**425 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5A80000000000000;

    #10 $display("\n2**424 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5A70000000000000;

    #10 $display("\n2**423 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5A60000000000000;

    #10 $display("\n2**422 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5A50000000000000;

    #10 $display("\n2**421 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5A40000000000000;

    #10 $display("\n2**420 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5A30000000000000;

    #10 $display("\n2**419 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5A20000000000000;

    #10 $display("\n2**418 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5A10000000000000;

    #10 $display("\n2**417 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5A00000000000000;

    #10 $display("\n2**416 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h59F0000000000000;

    #10 $display("\n2**415 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h59E0000000000000;

    #10 $display("\n2**414 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h59D0000000000000;

    #10 $display("\n2**413 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h59C0000000000000;

    #10 $display("\n2**412 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h59B0000000000000;

    #10 $display("\n2**411 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h59A0000000000000;

    #10 $display("\n2**410 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5990000000000000;

    #10 $display("\n2**409 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5980000000000000;

    #10 $display("\n2**408 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5970000000000000;

    #10 $display("\n2**407 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5960000000000000;

    #10 $display("\n2**406 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5950000000000000;

    #10 $display("\n2**405 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5940000000000000;

    #10 $display("\n2**404 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5930000000000000;

    #10 $display("\n2**403 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5920000000000000;

    #10 $display("\n2**402 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5910000000000000;

    #10 $display("\n2**401 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5900000000000000;

    #10 $display("\n2**400 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h58F0000000000000;

    #10 $display("\n2**399 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h58E0000000000000;

    #10 $display("\n2**398 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h58D0000000000000;

    #10 $display("\n2**397 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h58C0000000000000;

    #10 $display("\n2**396 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h58B0000000000000;

    #10 $display("\n2**395 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h58A0000000000000;

    #10 $display("\n2**394 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5890000000000000;

    #10 $display("\n2**393 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5880000000000000;

    #10 $display("\n2**392 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5870000000000000;

    #10 $display("\n2**391 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5860000000000000;

    #10 $display("\n2**390 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5850000000000000;

    #10 $display("\n2**389 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5840000000000000;

    #10 $display("\n2**388 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5830000000000000;

    #10 $display("\n2**387 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5820000000000000;

    #10 $display("\n2**386 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5810000000000000;

    #10 $display("\n2**385 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5800000000000000;

    #10 $display("\n2**384 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h57F0000000000000;

    #10 $display("\n2**383 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h57E0000000000000;

    #10 $display("\n2**382 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h57D0000000000000;

    #10 $display("\n2**381 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h57C0000000000000;

    #10 $display("\n2**380 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h57B0000000000000;

    #10 $display("\n2**379 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h57A0000000000000;

    #10 $display("\n2**378 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5790000000000000;

    #10 $display("\n2**377 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5780000000000000;

    #10 $display("\n2**376 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5770000000000000;

    #10 $display("\n2**375 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5760000000000000;

    #10 $display("\n2**374 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5750000000000000;

    #10 $display("\n2**373 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5740000000000000;

    #10 $display("\n2**372 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5730000000000000;

    #10 $display("\n2**371 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5720000000000000;

    #10 $display("\n2**370 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5710000000000000;

    #10 $display("\n2**369 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5700000000000000;

    #10 $display("\n2**368 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h56F0000000000000;

    #10 $display("\n2**367 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h56E0000000000000;

    #10 $display("\n2**366 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h56D0000000000000;

    #10 $display("\n2**365 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h56C0000000000000;

    #10 $display("\n2**364 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h56B0000000000000;

    #10 $display("\n2**363 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h56A0000000000000;

    #10 $display("\n2**362 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5690000000000000;

    #10 $display("\n2**361 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5680000000000000;

    #10 $display("\n2**360 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5670000000000000;

    #10 $display("\n2**359 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5660000000000000;

    #10 $display("\n2**358 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5650000000000000;

    #10 $display("\n2**357 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5640000000000000;

    #10 $display("\n2**356 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5630000000000000;

    #10 $display("\n2**355 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5620000000000000;

    #10 $display("\n2**354 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5610000000000000;

    #10 $display("\n2**353 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5600000000000000;

    #10 $display("\n2**352 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h55F0000000000000;

    #10 $display("\n2**351 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h55E0000000000000;

    #10 $display("\n2**350 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h55D0000000000000;

    #10 $display("\n2**349 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h55C0000000000000;

    #10 $display("\n2**348 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h55B0000000000000;

    #10 $display("\n2**347 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h55A0000000000000;

    #10 $display("\n2**346 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5590000000000000;

    #10 $display("\n2**345 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5580000000000000;

    #10 $display("\n2**344 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5570000000000000;

    #10 $display("\n2**343 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5560000000000000;

    #10 $display("\n2**342 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5550000000000000;

    #10 $display("\n2**341 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5540000000000000;

    #10 $display("\n2**340 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5530000000000000;

    #10 $display("\n2**339 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5520000000000000;

    #10 $display("\n2**338 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5510000000000000;

    #10 $display("\n2**337 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5500000000000000;

    #10 $display("\n2**336 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h54F0000000000000;

    #10 $display("\n2**335 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h54E0000000000000;

    #10 $display("\n2**334 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h54D0000000000000;

    #10 $display("\n2**333 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h54C0000000000000;

    #10 $display("\n2**332 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h54B0000000000000;

    #10 $display("\n2**331 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h54A0000000000000;

    #10 $display("\n2**330 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5490000000000000;

    #10 $display("\n2**329 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5480000000000000;

    #10 $display("\n2**328 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5470000000000000;

    #10 $display("\n2**327 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5460000000000000;

    #10 $display("\n2**326 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5450000000000000;

    #10 $display("\n2**325 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5440000000000000;

    #10 $display("\n2**324 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5430000000000000;

    #10 $display("\n2**323 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5420000000000000;

    #10 $display("\n2**322 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5410000000000000;

    #10 $display("\n2**321 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5400000000000000;

    #10 $display("\n2**320 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h53F0000000000000;

    #10 $display("\n2**319 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h53E0000000000000;

    #10 $display("\n2**318 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h53D0000000000000;

    #10 $display("\n2**317 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h53C0000000000000;

    #10 $display("\n2**316 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h53B0000000000000;

    #10 $display("\n2**315 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h53A0000000000000;

    #10 $display("\n2**314 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5390000000000000;

    #10 $display("\n2**313 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5380000000000000;

    #10 $display("\n2**312 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5370000000000000;

    #10 $display("\n2**311 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5360000000000000;

    #10 $display("\n2**310 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5350000000000000;

    #10 $display("\n2**309 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5340000000000000;

    #10 $display("\n2**308 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5330000000000000;

    #10 $display("\n2**307 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5320000000000000;

    #10 $display("\n2**306 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5310000000000000;

    #10 $display("\n2**305 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5300000000000000;

    #10 $display("\n2**304 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h52F0000000000000;

    #10 $display("\n2**303 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h52E0000000000000;

    #10 $display("\n2**302 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h52D0000000000000;

    #10 $display("\n2**301 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h52C0000000000000;

    #10 $display("\n2**300 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h52B0000000000000;

    #10 $display("\n2**299 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h52A0000000000000;

    #10 $display("\n2**298 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5290000000000000;

    #10 $display("\n2**297 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5280000000000000;

    #10 $display("\n2**296 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5270000000000000;

    #10 $display("\n2**295 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5260000000000000;

    #10 $display("\n2**294 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5250000000000000;

    #10 $display("\n2**293 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5240000000000000;

    #10 $display("\n2**292 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5230000000000000;

    #10 $display("\n2**291 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5220000000000000;

    #10 $display("\n2**290 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5210000000000000;

    #10 $display("\n2**289 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5200000000000000;

    #10 $display("\n2**288 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h51F0000000000000;

    #10 $display("\n2**287 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h51E0000000000000;

    #10 $display("\n2**286 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h51D0000000000000;

    #10 $display("\n2**285 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h51C0000000000000;

    #10 $display("\n2**284 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h51B0000000000000;

    #10 $display("\n2**283 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h51A0000000000000;

    #10 $display("\n2**282 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5190000000000000;

    #10 $display("\n2**281 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5180000000000000;

    #10 $display("\n2**280 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5170000000000000;

    #10 $display("\n2**279 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5160000000000000;

    #10 $display("\n2**278 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5150000000000000;

    #10 $display("\n2**277 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5140000000000000;

    #10 $display("\n2**276 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5130000000000000;

    #10 $display("\n2**275 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5120000000000000;

    #10 $display("\n2**274 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5110000000000000;

    #10 $display("\n2**273 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5100000000000000;

    #10 $display("\n2**272 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h50F0000000000000;

    #10 $display("\n2**271 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h50E0000000000000;

    #10 $display("\n2**270 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h50D0000000000000;

    #10 $display("\n2**269 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h50C0000000000000;

    #10 $display("\n2**268 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h50B0000000000000;

    #10 $display("\n2**267 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h50A0000000000000;

    #10 $display("\n2**266 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5090000000000000;

    #10 $display("\n2**265 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5080000000000000;

    #10 $display("\n2**264 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5070000000000000;

    #10 $display("\n2**263 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5060000000000000;

    #10 $display("\n2**262 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5050000000000000;

    #10 $display("\n2**261 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5040000000000000;

    #10 $display("\n2**260 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5030000000000000;

    #10 $display("\n2**259 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5020000000000000;

    #10 $display("\n2**258 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5010000000000000;

    #10 $display("\n2**257 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h5000000000000000;

    #10 $display("\n2**256 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4FF0000000000000;

    #10 $display("\n2**255 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4FE0000000000000;

    #10 $display("\n2**254 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4FD0000000000000;

    #10 $display("\n2**253 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4FC0000000000000;

    #10 $display("\n2**252 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4FB0000000000000;

    #10 $display("\n2**251 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4FA0000000000000;

    #10 $display("\n2**250 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4F90000000000000;

    #10 $display("\n2**249 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4F80000000000000;

    #10 $display("\n2**248 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4F70000000000000;

    #10 $display("\n2**247 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4F60000000000000;

    #10 $display("\n2**246 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4F50000000000000;

    #10 $display("\n2**245 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4F40000000000000;

    #10 $display("\n2**244 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4F30000000000000;

    #10 $display("\n2**243 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4F20000000000000;

    #10 $display("\n2**242 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4F10000000000000;

    #10 $display("\n2**241 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4F00000000000000;

    #10 $display("\n2**240 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4EF0000000000000;

    #10 $display("\n2**239 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4EE0000000000000;

    #10 $display("\n2**238 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4ED0000000000000;

    #10 $display("\n2**237 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4EC0000000000000;

    #10 $display("\n2**236 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4EB0000000000000;

    #10 $display("\n2**235 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4EA0000000000000;

    #10 $display("\n2**234 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4E90000000000000;

    #10 $display("\n2**233 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4E80000000000000;

    #10 $display("\n2**232 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4E70000000000000;

    #10 $display("\n2**231 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4E60000000000000;

    #10 $display("\n2**230 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4E50000000000000;

    #10 $display("\n2**229 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4E40000000000000;

    #10 $display("\n2**228 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4E30000000000000;

    #10 $display("\n2**227 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4E20000000000000;

    #10 $display("\n2**226 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4E10000000000000;

    #10 $display("\n2**225 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4E00000000000000;

    #10 $display("\n2**224 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4DF0000000000000;

    #10 $display("\n2**223 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4DE0000000000000;

    #10 $display("\n2**222 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4DD0000000000000;

    #10 $display("\n2**221 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4DC0000000000000;

    #10 $display("\n2**220 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4DB0000000000000;

    #10 $display("\n2**219 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4DA0000000000000;

    #10 $display("\n2**218 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4D90000000000000;

    #10 $display("\n2**217 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4D80000000000000;

    #10 $display("\n2**216 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4D70000000000000;

    #10 $display("\n2**215 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4D60000000000000;

    #10 $display("\n2**214 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4D50000000000000;

    #10 $display("\n2**213 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4D40000000000000;

    #10 $display("\n2**212 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4D30000000000000;

    #10 $display("\n2**211 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4D20000000000000;

    #10 $display("\n2**210 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4D10000000000000;

    #10 $display("\n2**209 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4D00000000000000;

    #10 $display("\n2**208 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4CF0000000000000;

    #10 $display("\n2**207 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4CE0000000000000;

    #10 $display("\n2**206 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4CD0000000000000;

    #10 $display("\n2**205 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4CC0000000000000;

    #10 $display("\n2**204 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4CB0000000000000;

    #10 $display("\n2**203 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4CA0000000000000;

    #10 $display("\n2**202 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4C90000000000000;

    #10 $display("\n2**201 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4C80000000000000;

    #10 $display("\n2**200 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4C70000000000000;

    #10 $display("\n2**199 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4C60000000000000;

    #10 $display("\n2**198 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4C50000000000000;

    #10 $display("\n2**197 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4C40000000000000;

    #10 $display("\n2**196 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4C30000000000000;

    #10 $display("\n2**195 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4C20000000000000;

    #10 $display("\n2**194 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4C10000000000000;

    #10 $display("\n2**193 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4C00000000000000;

    #10 $display("\n2**192 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4BF0000000000000;

    #10 $display("\n2**191 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4BE0000000000000;

    #10 $display("\n2**190 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4BD0000000000000;

    #10 $display("\n2**189 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4BC0000000000000;

    #10 $display("\n2**188 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4BB0000000000000;

    #10 $display("\n2**187 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4BA0000000000000;

    #10 $display("\n2**186 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4B90000000000000;

    #10 $display("\n2**185 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4B80000000000000;

    #10 $display("\n2**184 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4B70000000000000;

    #10 $display("\n2**183 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4B60000000000000;

    #10 $display("\n2**182 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4B50000000000000;

    #10 $display("\n2**181 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4B40000000000000;

    #10 $display("\n2**180 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4B30000000000000;

    #10 $display("\n2**179 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4B20000000000000;

    #10 $display("\n2**178 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4B10000000000000;

    #10 $display("\n2**177 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4B00000000000000;

    #10 $display("\n2**176 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4AF0000000000000;

    #10 $display("\n2**175 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4AE0000000000000;

    #10 $display("\n2**174 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4AD0000000000000;

    #10 $display("\n2**173 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4AC0000000000000;

    #10 $display("\n2**172 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4AB0000000000000;

    #10 $display("\n2**171 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4AA0000000000000;

    #10 $display("\n2**170 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4A90000000000000;

    #10 $display("\n2**169 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4A80000000000000;

    #10 $display("\n2**168 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4A70000000000000;

    #10 $display("\n2**167 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4A60000000000000;

    #10 $display("\n2**166 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4A50000000000000;

    #10 $display("\n2**165 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4A40000000000000;

    #10 $display("\n2**164 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4A30000000000000;

    #10 $display("\n2**163 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4A20000000000000;

    #10 $display("\n2**162 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4A10000000000000;

    #10 $display("\n2**161 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4A00000000000000;

    #10 $display("\n2**160 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h49F0000000000000;

    #10 $display("\n2**159 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h49E0000000000000;

    #10 $display("\n2**158 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h49D0000000000000;

    #10 $display("\n2**157 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h49C0000000000000;

    #10 $display("\n2**156 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h49B0000000000000;

    #10 $display("\n2**155 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h49A0000000000000;

    #10 $display("\n2**154 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4990000000000000;

    #10 $display("\n2**153 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4980000000000000;

    #10 $display("\n2**152 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4970000000000000;

    #10 $display("\n2**151 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4960000000000000;

    #10 $display("\n2**150 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4950000000000000;

    #10 $display("\n2**149 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4940000000000000;

    #10 $display("\n2**148 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4930000000000000;

    #10 $display("\n2**147 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4920000000000000;

    #10 $display("\n2**146 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4910000000000000;

    #10 $display("\n2**145 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4900000000000000;

    #10 $display("\n2**144 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h48F0000000000000;

    #10 $display("\n2**143 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h48E0000000000000;

    #10 $display("\n2**142 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h48D0000000000000;

    #10 $display("\n2**141 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h48C0000000000000;

    #10 $display("\n2**140 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h48B0000000000000;

    #10 $display("\n2**139 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h48A0000000000000;

    #10 $display("\n2**138 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4890000000000000;

    #10 $display("\n2**137 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4880000000000000;

    #10 $display("\n2**136 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4870000000000000;

    #10 $display("\n2**135 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4860000000000000;

    #10 $display("\n2**134 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4850000000000000;

    #10 $display("\n2**133 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4840000000000000;

    #10 $display("\n2**132 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4830000000000000;

    #10 $display("\n2**131 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4820000000000000;

    #10 $display("\n2**130 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4810000000000000;

    #10 $display("\n2**129 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4800000000000000;

    #10 $display("\n2**128 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h47F0000000000000;

    #10 $display("\n2**127 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h47E0000000000000;

    #10 $display("\n2**126 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h47D0000000000000;

    #10 $display("\n2**125 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h47C0000000000000;

    #10 $display("\n2**124 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h47B0000000000000;

    #10 $display("\n2**123 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h47A0000000000000;

    #10 $display("\n2**122 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4790000000000000;

    #10 $display("\n2**121 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4780000000000000;

    #10 $display("\n2**120 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4770000000000000;

    #10 $display("\n2**119 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4760000000000000;

    #10 $display("\n2**118 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4750000000000000;

    #10 $display("\n2**117 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4740000000000000;

    #10 $display("\n2**116 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4730000000000000;

    #10 $display("\n2**115 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4720000000000000;

    #10 $display("\n2**114 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4710000000000000;

    #10 $display("\n2**113 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4700000000000000;

    #10 $display("\n2**112 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h46F0000000000000;

    #10 $display("\n2**111 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h46E0000000000000;

    #10 $display("\n2**110 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h46D0000000000000;

    #10 $display("\n2**109 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h46C0000000000000;

    #10 $display("\n2**108 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h46B0000000000000;

    #10 $display("\n2**107 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h46A0000000000000;

    #10 $display("\n2**106 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4690000000000000;

    #10 $display("\n2**105 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4680000000000000;

    #10 $display("\n2**104 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4670000000000000;

    #10 $display("\n2**103 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4660000000000000;

    #10 $display("\n2**102 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4650000000000000;

    #10 $display("\n2**101 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4640000000000000;

    #10 $display("\n2**100 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4630000000000000;

    #10 $display("\n2**99 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4620000000000000;

    #10 $display("\n2**98 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4610000000000000;

    #10 $display("\n2**97 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4600000000000000;

    #10 $display("\n2**96 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h45F0000000000000;

    #10 $display("\n2**95 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h45E0000000000000;

    #10 $display("\n2**94 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h45D0000000000000;

    #10 $display("\n2**93 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h45C0000000000000;

    #10 $display("\n2**92 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h45B0000000000000;

    #10 $display("\n2**91 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h45A0000000000000;

    #10 $display("\n2**90 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4590000000000000;

    #10 $display("\n2**89 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4580000000000000;

    #10 $display("\n2**88 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4570000000000000;

    #10 $display("\n2**87 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4560000000000000;

    #10 $display("\n2**86 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4550000000000000;

    #10 $display("\n2**85 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4540000000000000;

    #10 $display("\n2**84 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4530000000000000;

    #10 $display("\n2**83 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4520000000000000;

    #10 $display("\n2**82 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4510000000000000;

    #10 $display("\n2**81 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4500000000000000;

    #10 $display("\n2**80 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h44F0000000000000;

    #10 $display("\n2**79 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h44E0000000000000;

    #10 $display("\n2**78 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h44D0000000000000;

    #10 $display("\n2**77 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h44C0000000000000;

    #10 $display("\n2**76 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h44B0000000000000;

    #10 $display("\n2**75 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h44A0000000000000;

    #10 $display("\n2**74 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4490000000000000;

    #10 $display("\n2**73 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4480000000000000;

    #10 $display("\n2**72 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4470000000000000;

    #10 $display("\n2**71 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4460000000000000;

    #10 $display("\n2**70 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4450000000000000;

    #10 $display("\n2**69 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4440000000000000;

    #10 $display("\n2**68 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4430000000000000;

    #10 $display("\n2**67 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4420000000000000;

    #10 $display("\n2**66 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4410000000000000;

    #10 $display("\n2**65 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4400000000000000;

    #10 $display("\n2**64 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h43F0000000000000;

    #10 $display("\n2**63 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h43E0000000000000;

    #10 $display("\n2**62 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h43D0000000000000;

    #10 $display("\n2**61 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h43C0000000000000;

    #10 $display("\n2**60 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h43B0000000000000;

    #10 $display("\n2**59 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h43A0000000000000;

    #10 $display("\n2**58 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4390000000000000;

    #10 $display("\n2**57 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4380000000000000;

    #10 $display("\n2**56 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4370000000000000;

    #10 $display("\n2**55 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4360000000000000;

    #10 $display("\n2**54 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4350000000000000;

    #10 $display("\n2**53 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4340000000000000;

    #10 $display("\n2**52 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4330000000000000;

    #10 $display("\n2**51 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4320000000000000;

    #10 $display("\n2**50 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4310000000000000;

    #10 $display("\n2**49 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4300000000000000;

    #10 $display("\n2**48 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h42F0000000000000;

    #10 $display("\n2**47 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h42E0000000000000;

    #10 $display("\n2**46 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h42D0000000000000;

    #10 $display("\n2**45 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h42C0000000000000;

    #10 $display("\n2**44 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h42B0000000000000;

    #10 $display("\n2**43 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h42A0000000000000;

    #10 $display("\n2**42 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4290000000000000;

    #10 $display("\n2**41 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4280000000000000;

    #10 $display("\n2**40 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4270000000000000;

    #10 $display("\n2**39 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4260000000000000;

    #10 $display("\n2**38 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4250000000000000;

    #10 $display("\n2**37 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4240000000000000;

    #10 $display("\n2**36 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4230000000000000;

    #10 $display("\n2**35 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4220000000000000;

    #10 $display("\n2**34 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4210000000000000;

    #10 $display("\n2**33 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4200000000000000;

    #10 $display("\n2**32 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h41F0000000000000;

    #10 $display("\n2**31 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h41E0000000000000;

    #10 $display("\n2**30 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h41D0000000000000;

    #10 $display("\n2**29 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h41C0000000000000;

    #10 $display("\n2**28 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h41B0000000000000;

    #10 $display("\n2**27 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h41A0000000000000;

    #10 $display("\n2**26 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4190000000000000;

    #10 $display("\n2**25 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4180000000000000;

    #10 $display("\n2**24 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4170000000000000;

    #10 $display("\n2**23 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4160000000000000;

    #10 $display("\n2**22 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4150000000000000;

    #10 $display("\n2**21 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4140000000000000;

    #10 $display("\n2**20 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4130000000000000;

    #10 $display("\n2**19 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4120000000000000;

    #10 $display("\n2**18 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4110000000000000;

    #10 $display("\n2**17 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4100000000000000;

    #10 $display("\n2**16 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h40F0000000000000;

    #10 $display("\n2**15 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h40E0000000000000;

    #10 $display("\n2**14 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h40D0000000000000;

    #10 $display("\n2**13 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h40C0000000000000;

    #10 $display("\n2**12 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h40B0000000000000;

    #10 $display("\n2**11 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h40A0000000000000;

    #10 $display("\n2**10 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4090000000000000;

    #10 $display("\n2**9 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4080000000000000;

    #10 $display("\n2**8 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4070000000000000;

    #10 $display("\n2**7 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4060000000000000;

    #10 $display("\n2**6 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4050000000000000;

    #10 $display("\n2**5 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4040000000000000;

    #10 $display("\n2**4 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4030000000000000;

    #10 $display("\n2**3 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4020000000000000;

    #10 $display("\n2**2 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4010000000000000;

    #10 $display("\n2**1 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h4000000000000000;

    #10 $display("\n2**0 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3FF0000000000000;

    #10 $display("\n2**-1 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3FE0000000000000;

    #10 $display("\n2**-2 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3FD0000000000000;

    #10 $display("\n2**-3 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3FC0000000000000;

    #10 $display("\n2**-4 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3FB0000000000000;

    #10 $display("\n2**-5 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3FA0000000000000;

    #10 $display("\n2**-6 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3F90000000000000;

    #10 $display("\n2**-7 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3F80000000000000;

    #10 $display("\n2**-8 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3F70000000000000;

    #10 $display("\n2**-9 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3F60000000000000;

    #10 $display("\n2**-10 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3F50000000000000;

    #10 $display("\n2**-11 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3F40000000000000;

    #10 $display("\n2**-12 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3F30000000000000;

    #10 $display("\n2**-13 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3F20000000000000;

    #10 $display("\n2**-14 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3F10000000000000;

    #10 $display("\n2**-15 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3F00000000000000;

    #10 $display("\n2**-16 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3EF0000000000000;

    #10 $display("\n2**-17 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3EE0000000000000;

    #10 $display("\n2**-18 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3ED0000000000000;

    #10 $display("\n2**-19 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3EC0000000000000;

    #10 $display("\n2**-20 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3EB0000000000000;

    #10 $display("\n2**-21 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3EA0000000000000;

    #10 $display("\n2**-22 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3E90000000000000;

    #10 $display("\n2**-23 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3E80000000000000;

    #10 $display("\n2**-24 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3E70000000000000;

    #10 $display("\n2**-25 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3E60000000000000;

    #10 $display("\n2**-26 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3E50000000000000;

    #10 $display("\n2**-27 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3E40000000000000;

    #10 $display("\n2**-28 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3E30000000000000;

    #10 $display("\n2**-29 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3E20000000000000;

    #10 $display("\n2**-30 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3E10000000000000;

    #10 $display("\n2**-31 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3E00000000000000;

    #10 $display("\n2**-32 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3DF0000000000000;

    #10 $display("\n2**-33 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3DE0000000000000;

    #10 $display("\n2**-34 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3DD0000000000000;

    #10 $display("\n2**-35 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3DC0000000000000;

    #10 $display("\n2**-36 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3DB0000000000000;

    #10 $display("\n2**-37 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3DA0000000000000;

    #10 $display("\n2**-38 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3D90000000000000;

    #10 $display("\n2**-39 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3D80000000000000;

    #10 $display("\n2**-40 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3D70000000000000;

    #10 $display("\n2**-41 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3D60000000000000;

    #10 $display("\n2**-42 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3D50000000000000;

    #10 $display("\n2**-43 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3D40000000000000;

    #10 $display("\n2**-44 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3D30000000000000;

    #10 $display("\n2**-45 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3D20000000000000;

    #10 $display("\n2**-46 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3D10000000000000;

    #10 $display("\n2**-47 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3D00000000000000;

    #10 $display("\n2**-48 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3CF0000000000000;

    #10 $display("\n2**-49 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3CE0000000000000;

    #10 $display("\n2**-50 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3CD0000000000000;

    #10 $display("\n2**-51 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3CC0000000000000;

    #10 $display("\n2**-52 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3CB0000000000000;

    #10 $display("\n2**-53 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3CA0000000000000;

    #10 $display("\n2**-54 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3C90000000000000;

    #10 $display("\n2**-55 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3C80000000000000;

    #10 $display("\n2**-56 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3C70000000000000;

    #10 $display("\n2**-57 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3C60000000000000;

    #10 $display("\n2**-58 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3C50000000000000;

    #10 $display("\n2**-59 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3C40000000000000;

    #10 $display("\n2**-60 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3C30000000000000;

    #10 $display("\n2**-61 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3C20000000000000;

    #10 $display("\n2**-62 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3C10000000000000;

    #10 $display("\n2**-63 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3C00000000000000;

    #10 $display("\n2**-64 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3BF0000000000000;

    #10 $display("\n2**-65 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3BE0000000000000;

    #10 $display("\n2**-66 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3BD0000000000000;

    #10 $display("\n2**-67 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3BC0000000000000;

    #10 $display("\n2**-68 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3BB0000000000000;

    #10 $display("\n2**-69 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3BA0000000000000;

    #10 $display("\n2**-70 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3B90000000000000;

    #10 $display("\n2**-71 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3B80000000000000;

    #10 $display("\n2**-72 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3B70000000000000;

    #10 $display("\n2**-73 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3B60000000000000;

    #10 $display("\n2**-74 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3B50000000000000;

    #10 $display("\n2**-75 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3B40000000000000;

    #10 $display("\n2**-76 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3B30000000000000;

    #10 $display("\n2**-77 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3B20000000000000;

    #10 $display("\n2**-78 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3B10000000000000;

    #10 $display("\n2**-79 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3B00000000000000;

    #10 $display("\n2**-80 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3AF0000000000000;

    #10 $display("\n2**-81 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3AE0000000000000;

    #10 $display("\n2**-82 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3AD0000000000000;

    #10 $display("\n2**-83 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3AC0000000000000;

    #10 $display("\n2**-84 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3AB0000000000000;

    #10 $display("\n2**-85 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3AA0000000000000;

    #10 $display("\n2**-86 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3A90000000000000;

    #10 $display("\n2**-87 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3A80000000000000;

    #10 $display("\n2**-88 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3A70000000000000;

    #10 $display("\n2**-89 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3A60000000000000;

    #10 $display("\n2**-90 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3A50000000000000;

    #10 $display("\n2**-91 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3A40000000000000;

    #10 $display("\n2**-92 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3A30000000000000;

    #10 $display("\n2**-93 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3A20000000000000;

    #10 $display("\n2**-94 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3A10000000000000;

    #10 $display("\n2**-95 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3A00000000000000;

    #10 $display("\n2**-96 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h39F0000000000000;

    #10 $display("\n2**-97 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h39E0000000000000;

    #10 $display("\n2**-98 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h39D0000000000000;

    #10 $display("\n2**-99 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h39C0000000000000;

    #10 $display("\n2**-100 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h39B0000000000000;

    #10 $display("\n2**-101 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h39A0000000000000;

    #10 $display("\n2**-102 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3990000000000000;

    #10 $display("\n2**-103 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3980000000000000;

    #10 $display("\n2**-104 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3970000000000000;

    #10 $display("\n2**-105 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3960000000000000;

    #10 $display("\n2**-106 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3950000000000000;

    #10 $display("\n2**-107 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3940000000000000;

    #10 $display("\n2**-108 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3930000000000000;

    #10 $display("\n2**-109 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3920000000000000;

    #10 $display("\n2**-110 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3910000000000000;

    #10 $display("\n2**-111 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3900000000000000;

    #10 $display("\n2**-112 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h38F0000000000000;

    #10 $display("\n2**-113 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h38E0000000000000;

    #10 $display("\n2**-114 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h38D0000000000000;

    #10 $display("\n2**-115 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h38C0000000000000;

    #10 $display("\n2**-116 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h38B0000000000000;

    #10 $display("\n2**-117 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h38A0000000000000;

    #10 $display("\n2**-118 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3890000000000000;

    #10 $display("\n2**-119 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3880000000000000;

    #10 $display("\n2**-120 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3870000000000000;

    #10 $display("\n2**-121 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3860000000000000;

    #10 $display("\n2**-122 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3850000000000000;

    #10 $display("\n2**-123 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3840000000000000;

    #10 $display("\n2**-124 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3830000000000000;

    #10 $display("\n2**-125 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3820000000000000;

    #10 $display("\n2**-126 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3810000000000000;

    #10 $display("\n2**-127 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3800000000000000;

    #10 $display("\n2**-128 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h37F0000000000000;

    #10 $display("\n2**-129 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h37E0000000000000;

    #10 $display("\n2**-130 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h37D0000000000000;

    #10 $display("\n2**-131 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h37C0000000000000;

    #10 $display("\n2**-132 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h37B0000000000000;

    #10 $display("\n2**-133 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h37A0000000000000;

    #10 $display("\n2**-134 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3790000000000000;

    #10 $display("\n2**-135 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3780000000000000;

    #10 $display("\n2**-136 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3770000000000000;

    #10 $display("\n2**-137 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3760000000000000;

    #10 $display("\n2**-138 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3750000000000000;

    #10 $display("\n2**-139 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3740000000000000;

    #10 $display("\n2**-140 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3730000000000000;

    #10 $display("\n2**-141 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3720000000000000;

    #10 $display("\n2**-142 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3710000000000000;

    #10 $display("\n2**-143 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3700000000000000;

    #10 $display("\n2**-144 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h36F0000000000000;

    #10 $display("\n2**-145 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h36E0000000000000;

    #10 $display("\n2**-146 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h36D0000000000000;

    #10 $display("\n2**-147 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h36C0000000000000;

    #10 $display("\n2**-148 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h36B0000000000000;

    #10 $display("\n2**-149 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h36A0000000000000;

    #10 $display("\n2**-150 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3690000000000000;

    #10 $display("\n2**-151 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3680000000000000;

    #10 $display("\n2**-152 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3670000000000000;

    #10 $display("\n2**-153 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3660000000000000;

    #10 $display("\n2**-154 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3650000000000000;

    #10 $display("\n2**-155 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3640000000000000;

    #10 $display("\n2**-156 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3630000000000000;

    #10 $display("\n2**-157 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3620000000000000;

    #10 $display("\n2**-158 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3610000000000000;

    #10 $display("\n2**-159 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3600000000000000;

    #10 $display("\n2**-160 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h35F0000000000000;

    #10 $display("\n2**-161 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h35E0000000000000;

    #10 $display("\n2**-162 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h35D0000000000000;

    #10 $display("\n2**-163 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h35C0000000000000;

    #10 $display("\n2**-164 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h35B0000000000000;

    #10 $display("\n2**-165 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h35A0000000000000;

    #10 $display("\n2**-166 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3590000000000000;

    #10 $display("\n2**-167 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3580000000000000;

    #10 $display("\n2**-168 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3570000000000000;

    #10 $display("\n2**-169 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3560000000000000;

    #10 $display("\n2**-170 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3550000000000000;

    #10 $display("\n2**-171 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3540000000000000;

    #10 $display("\n2**-172 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3530000000000000;

    #10 $display("\n2**-173 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3520000000000000;

    #10 $display("\n2**-174 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3510000000000000;

    #10 $display("\n2**-175 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3500000000000000;

    #10 $display("\n2**-176 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h34F0000000000000;

    #10 $display("\n2**-177 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h34E0000000000000;

    #10 $display("\n2**-178 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h34D0000000000000;

    #10 $display("\n2**-179 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h34C0000000000000;

    #10 $display("\n2**-180 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h34B0000000000000;

    #10 $display("\n2**-181 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h34A0000000000000;

    #10 $display("\n2**-182 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3490000000000000;

    #10 $display("\n2**-183 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3480000000000000;

    #10 $display("\n2**-184 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3470000000000000;

    #10 $display("\n2**-185 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3460000000000000;

    #10 $display("\n2**-186 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3450000000000000;

    #10 $display("\n2**-187 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3440000000000000;

    #10 $display("\n2**-188 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3430000000000000;

    #10 $display("\n2**-189 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3420000000000000;

    #10 $display("\n2**-190 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3410000000000000;

    #10 $display("\n2**-191 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3400000000000000;

    #10 $display("\n2**-192 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h33F0000000000000;

    #10 $display("\n2**-193 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h33E0000000000000;

    #10 $display("\n2**-194 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h33D0000000000000;

    #10 $display("\n2**-195 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h33C0000000000000;

    #10 $display("\n2**-196 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h33B0000000000000;

    #10 $display("\n2**-197 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h33A0000000000000;

    #10 $display("\n2**-198 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3390000000000000;

    #10 $display("\n2**-199 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3380000000000000;

    #10 $display("\n2**-200 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3370000000000000;

    #10 $display("\n2**-201 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3360000000000000;

    #10 $display("\n2**-202 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3350000000000000;

    #10 $display("\n2**-203 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3340000000000000;

    #10 $display("\n2**-204 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3330000000000000;

    #10 $display("\n2**-205 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3320000000000000;

    #10 $display("\n2**-206 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3310000000000000;

    #10 $display("\n2**-207 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3300000000000000;

    #10 $display("\n2**-208 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h32F0000000000000;

    #10 $display("\n2**-209 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h32E0000000000000;

    #10 $display("\n2**-210 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h32D0000000000000;

    #10 $display("\n2**-211 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h32C0000000000000;

    #10 $display("\n2**-212 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h32B0000000000000;

    #10 $display("\n2**-213 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h32A0000000000000;

    #10 $display("\n2**-214 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3290000000000000;

    #10 $display("\n2**-215 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3280000000000000;

    #10 $display("\n2**-216 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3270000000000000;

    #10 $display("\n2**-217 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3260000000000000;

    #10 $display("\n2**-218 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3250000000000000;

    #10 $display("\n2**-219 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3240000000000000;

    #10 $display("\n2**-220 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3230000000000000;

    #10 $display("\n2**-221 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3220000000000000;

    #10 $display("\n2**-222 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3210000000000000;

    #10 $display("\n2**-223 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3200000000000000;

    #10 $display("\n2**-224 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h31F0000000000000;

    #10 $display("\n2**-225 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h31E0000000000000;

    #10 $display("\n2**-226 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h31D0000000000000;

    #10 $display("\n2**-227 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h31C0000000000000;

    #10 $display("\n2**-228 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h31B0000000000000;

    #10 $display("\n2**-229 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h31A0000000000000;

    #10 $display("\n2**-230 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3190000000000000;

    #10 $display("\n2**-231 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3180000000000000;

    #10 $display("\n2**-232 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3170000000000000;

    #10 $display("\n2**-233 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3160000000000000;

    #10 $display("\n2**-234 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3150000000000000;

    #10 $display("\n2**-235 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3140000000000000;

    #10 $display("\n2**-236 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3130000000000000;

    #10 $display("\n2**-237 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3120000000000000;

    #10 $display("\n2**-238 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3110000000000000;

    #10 $display("\n2**-239 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3100000000000000;

    #10 $display("\n2**-240 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h30F0000000000000;

    #10 $display("\n2**-241 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h30E0000000000000;

    #10 $display("\n2**-242 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h30D0000000000000;

    #10 $display("\n2**-243 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h30C0000000000000;

    #10 $display("\n2**-244 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h30B0000000000000;

    #10 $display("\n2**-245 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h30A0000000000000;

    #10 $display("\n2**-246 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3090000000000000;

    #10 $display("\n2**-247 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3080000000000000;

    #10 $display("\n2**-248 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3070000000000000;

    #10 $display("\n2**-249 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3060000000000000;

    #10 $display("\n2**-250 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3050000000000000;

    #10 $display("\n2**-251 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3040000000000000;

    #10 $display("\n2**-252 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3030000000000000;

    #10 $display("\n2**-253 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3020000000000000;

    #10 $display("\n2**-254 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3010000000000000;

    #10 $display("\n2**-255 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h3000000000000000;

    #10 $display("\n2**-256 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2FF0000000000000;

    #10 $display("\n2**-257 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2FE0000000000000;

    #10 $display("\n2**-258 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2FD0000000000000;

    #10 $display("\n2**-259 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2FC0000000000000;

    #10 $display("\n2**-260 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2FB0000000000000;

    #10 $display("\n2**-261 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2FA0000000000000;

    #10 $display("\n2**-262 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2F90000000000000;

    #10 $display("\n2**-263 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2F80000000000000;

    #10 $display("\n2**-264 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2F70000000000000;

    #10 $display("\n2**-265 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2F60000000000000;

    #10 $display("\n2**-266 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2F50000000000000;

    #10 $display("\n2**-267 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2F40000000000000;

    #10 $display("\n2**-268 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2F30000000000000;

    #10 $display("\n2**-269 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2F20000000000000;

    #10 $display("\n2**-270 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2F10000000000000;

    #10 $display("\n2**-271 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2F00000000000000;

    #10 $display("\n2**-272 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2EF0000000000000;

    #10 $display("\n2**-273 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2EE0000000000000;

    #10 $display("\n2**-274 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2ED0000000000000;

    #10 $display("\n2**-275 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2EC0000000000000;

    #10 $display("\n2**-276 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2EB0000000000000;

    #10 $display("\n2**-277 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2EA0000000000000;

    #10 $display("\n2**-278 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2E90000000000000;

    #10 $display("\n2**-279 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2E80000000000000;

    #10 $display("\n2**-280 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2E70000000000000;

    #10 $display("\n2**-281 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2E60000000000000;

    #10 $display("\n2**-282 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2E50000000000000;

    #10 $display("\n2**-283 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2E40000000000000;

    #10 $display("\n2**-284 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2E30000000000000;

    #10 $display("\n2**-285 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2E20000000000000;

    #10 $display("\n2**-286 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2E10000000000000;

    #10 $display("\n2**-287 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2E00000000000000;

    #10 $display("\n2**-288 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2DF0000000000000;

    #10 $display("\n2**-289 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2DE0000000000000;

    #10 $display("\n2**-290 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2DD0000000000000;

    #10 $display("\n2**-291 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2DC0000000000000;

    #10 $display("\n2**-292 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2DB0000000000000;

    #10 $display("\n2**-293 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2DA0000000000000;

    #10 $display("\n2**-294 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2D90000000000000;

    #10 $display("\n2**-295 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2D80000000000000;

    #10 $display("\n2**-296 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2D70000000000000;

    #10 $display("\n2**-297 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2D60000000000000;

    #10 $display("\n2**-298 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2D50000000000000;

    #10 $display("\n2**-299 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2D40000000000000;

    #10 $display("\n2**-300 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2D30000000000000;

    #10 $display("\n2**-301 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2D20000000000000;

    #10 $display("\n2**-302 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2D10000000000000;

    #10 $display("\n2**-303 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2D00000000000000;

    #10 $display("\n2**-304 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2CF0000000000000;

    #10 $display("\n2**-305 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2CE0000000000000;

    #10 $display("\n2**-306 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2CD0000000000000;

    #10 $display("\n2**-307 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2CC0000000000000;

    #10 $display("\n2**-308 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2CB0000000000000;

    #10 $display("\n2**-309 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2CA0000000000000;

    #10 $display("\n2**-310 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2C90000000000000;

    #10 $display("\n2**-311 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2C80000000000000;

    #10 $display("\n2**-312 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2C70000000000000;

    #10 $display("\n2**-313 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2C60000000000000;

    #10 $display("\n2**-314 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2C50000000000000;

    #10 $display("\n2**-315 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2C40000000000000;

    #10 $display("\n2**-316 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2C30000000000000;

    #10 $display("\n2**-317 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2C20000000000000;

    #10 $display("\n2**-318 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2C10000000000000;

    #10 $display("\n2**-319 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2C00000000000000;

    #10 $display("\n2**-320 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2BF0000000000000;

    #10 $display("\n2**-321 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2BE0000000000000;

    #10 $display("\n2**-322 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2BD0000000000000;

    #10 $display("\n2**-323 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2BC0000000000000;

    #10 $display("\n2**-324 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2BB0000000000000;

    #10 $display("\n2**-325 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2BA0000000000000;

    #10 $display("\n2**-326 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2B90000000000000;

    #10 $display("\n2**-327 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2B80000000000000;

    #10 $display("\n2**-328 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2B70000000000000;

    #10 $display("\n2**-329 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2B60000000000000;

    #10 $display("\n2**-330 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2B50000000000000;

    #10 $display("\n2**-331 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2B40000000000000;

    #10 $display("\n2**-332 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2B30000000000000;

    #10 $display("\n2**-333 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2B20000000000000;

    #10 $display("\n2**-334 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2B10000000000000;

    #10 $display("\n2**-335 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2B00000000000000;

    #10 $display("\n2**-336 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2AF0000000000000;

    #10 $display("\n2**-337 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2AE0000000000000;

    #10 $display("\n2**-338 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2AD0000000000000;

    #10 $display("\n2**-339 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2AC0000000000000;

    #10 $display("\n2**-340 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2AB0000000000000;

    #10 $display("\n2**-341 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2AA0000000000000;

    #10 $display("\n2**-342 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2A90000000000000;

    #10 $display("\n2**-343 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2A80000000000000;

    #10 $display("\n2**-344 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2A70000000000000;

    #10 $display("\n2**-345 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2A60000000000000;

    #10 $display("\n2**-346 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2A50000000000000;

    #10 $display("\n2**-347 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2A40000000000000;

    #10 $display("\n2**-348 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2A30000000000000;

    #10 $display("\n2**-349 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2A20000000000000;

    #10 $display("\n2**-350 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2A10000000000000;

    #10 $display("\n2**-351 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2A00000000000000;

    #10 $display("\n2**-352 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h29F0000000000000;

    #10 $display("\n2**-353 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h29E0000000000000;

    #10 $display("\n2**-354 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h29D0000000000000;

    #10 $display("\n2**-355 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h29C0000000000000;

    #10 $display("\n2**-356 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h29B0000000000000;

    #10 $display("\n2**-357 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h29A0000000000000;

    #10 $display("\n2**-358 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2990000000000000;

    #10 $display("\n2**-359 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2980000000000000;

    #10 $display("\n2**-360 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2970000000000000;

    #10 $display("\n2**-361 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2960000000000000;

    #10 $display("\n2**-362 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2950000000000000;

    #10 $display("\n2**-363 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2940000000000000;

    #10 $display("\n2**-364 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2930000000000000;

    #10 $display("\n2**-365 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2920000000000000;

    #10 $display("\n2**-366 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2910000000000000;

    #10 $display("\n2**-367 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2900000000000000;

    #10 $display("\n2**-368 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h28F0000000000000;

    #10 $display("\n2**-369 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h28E0000000000000;

    #10 $display("\n2**-370 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h28D0000000000000;

    #10 $display("\n2**-371 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h28C0000000000000;

    #10 $display("\n2**-372 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h28B0000000000000;

    #10 $display("\n2**-373 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h28A0000000000000;

    #10 $display("\n2**-374 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2890000000000000;

    #10 $display("\n2**-375 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2880000000000000;

    #10 $display("\n2**-376 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2870000000000000;

    #10 $display("\n2**-377 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2860000000000000;

    #10 $display("\n2**-378 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2850000000000000;

    #10 $display("\n2**-379 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2840000000000000;

    #10 $display("\n2**-380 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2830000000000000;

    #10 $display("\n2**-381 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2820000000000000;

    #10 $display("\n2**-382 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2810000000000000;

    #10 $display("\n2**-383 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2800000000000000;

    #10 $display("\n2**-384 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h27F0000000000000;

    #10 $display("\n2**-385 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h27E0000000000000;

    #10 $display("\n2**-386 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h27D0000000000000;

    #10 $display("\n2**-387 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h27C0000000000000;

    #10 $display("\n2**-388 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h27B0000000000000;

    #10 $display("\n2**-389 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h27A0000000000000;

    #10 $display("\n2**-390 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2790000000000000;

    #10 $display("\n2**-391 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2780000000000000;

    #10 $display("\n2**-392 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2770000000000000;

    #10 $display("\n2**-393 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2760000000000000;

    #10 $display("\n2**-394 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2750000000000000;

    #10 $display("\n2**-395 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2740000000000000;

    #10 $display("\n2**-396 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2730000000000000;

    #10 $display("\n2**-397 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2720000000000000;

    #10 $display("\n2**-398 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2710000000000000;

    #10 $display("\n2**-399 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2700000000000000;

    #10 $display("\n2**-400 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h26F0000000000000;

    #10 $display("\n2**-401 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h26E0000000000000;

    #10 $display("\n2**-402 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h26D0000000000000;

    #10 $display("\n2**-403 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h26C0000000000000;

    #10 $display("\n2**-404 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h26B0000000000000;

    #10 $display("\n2**-405 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h26A0000000000000;

    #10 $display("\n2**-406 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2690000000000000;

    #10 $display("\n2**-407 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2680000000000000;

    #10 $display("\n2**-408 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2670000000000000;

    #10 $display("\n2**-409 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2660000000000000;

    #10 $display("\n2**-410 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2650000000000000;

    #10 $display("\n2**-411 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2640000000000000;

    #10 $display("\n2**-412 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2630000000000000;

    #10 $display("\n2**-413 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2620000000000000;

    #10 $display("\n2**-414 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2610000000000000;

    #10 $display("\n2**-415 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2600000000000000;

    #10 $display("\n2**-416 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h25F0000000000000;

    #10 $display("\n2**-417 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h25E0000000000000;

    #10 $display("\n2**-418 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h25D0000000000000;

    #10 $display("\n2**-419 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h25C0000000000000;

    #10 $display("\n2**-420 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h25B0000000000000;

    #10 $display("\n2**-421 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h25A0000000000000;

    #10 $display("\n2**-422 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2590000000000000;

    #10 $display("\n2**-423 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2580000000000000;

    #10 $display("\n2**-424 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2570000000000000;

    #10 $display("\n2**-425 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2560000000000000;

    #10 $display("\n2**-426 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2550000000000000;

    #10 $display("\n2**-427 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2540000000000000;

    #10 $display("\n2**-428 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2530000000000000;

    #10 $display("\n2**-429 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2520000000000000;

    #10 $display("\n2**-430 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2510000000000000;

    #10 $display("\n2**-431 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2500000000000000;

    #10 $display("\n2**-432 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h24F0000000000000;

    #10 $display("\n2**-433 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h24E0000000000000;

    #10 $display("\n2**-434 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h24D0000000000000;

    #10 $display("\n2**-435 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h24C0000000000000;

    #10 $display("\n2**-436 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h24B0000000000000;

    #10 $display("\n2**-437 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h24A0000000000000;

    #10 $display("\n2**-438 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2490000000000000;

    #10 $display("\n2**-439 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2480000000000000;

    #10 $display("\n2**-440 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2470000000000000;

    #10 $display("\n2**-441 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2460000000000000;

    #10 $display("\n2**-442 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2450000000000000;

    #10 $display("\n2**-443 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2440000000000000;

    #10 $display("\n2**-444 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2430000000000000;

    #10 $display("\n2**-445 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2420000000000000;

    #10 $display("\n2**-446 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2410000000000000;

    #10 $display("\n2**-447 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2400000000000000;

    #10 $display("\n2**-448 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h23F0000000000000;

    #10 $display("\n2**-449 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h23E0000000000000;

    #10 $display("\n2**-450 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h23D0000000000000;

    #10 $display("\n2**-451 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h23C0000000000000;

    #10 $display("\n2**-452 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h23B0000000000000;

    #10 $display("\n2**-453 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h23A0000000000000;

    #10 $display("\n2**-454 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2390000000000000;

    #10 $display("\n2**-455 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2380000000000000;

    #10 $display("\n2**-456 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2370000000000000;

    #10 $display("\n2**-457 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2360000000000000;

    #10 $display("\n2**-458 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2350000000000000;

    #10 $display("\n2**-459 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2340000000000000;

    #10 $display("\n2**-460 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2330000000000000;

    #10 $display("\n2**-461 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2320000000000000;

    #10 $display("\n2**-462 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2310000000000000;

    #10 $display("\n2**-463 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2300000000000000;

    #10 $display("\n2**-464 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h22F0000000000000;

    #10 $display("\n2**-465 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h22E0000000000000;

    #10 $display("\n2**-466 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h22D0000000000000;

    #10 $display("\n2**-467 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h22C0000000000000;

    #10 $display("\n2**-468 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h22B0000000000000;

    #10 $display("\n2**-469 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h22A0000000000000;

    #10 $display("\n2**-470 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2290000000000000;

    #10 $display("\n2**-471 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2280000000000000;

    #10 $display("\n2**-472 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2270000000000000;

    #10 $display("\n2**-473 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2260000000000000;

    #10 $display("\n2**-474 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2250000000000000;

    #10 $display("\n2**-475 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2240000000000000;

    #10 $display("\n2**-476 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2230000000000000;

    #10 $display("\n2**-477 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2220000000000000;

    #10 $display("\n2**-478 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2210000000000000;

    #10 $display("\n2**-479 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2200000000000000;

    #10 $display("\n2**-480 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h21F0000000000000;

    #10 $display("\n2**-481 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h21E0000000000000;

    #10 $display("\n2**-482 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h21D0000000000000;

    #10 $display("\n2**-483 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h21C0000000000000;

    #10 $display("\n2**-484 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h21B0000000000000;

    #10 $display("\n2**-485 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h21A0000000000000;

    #10 $display("\n2**-486 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2190000000000000;

    #10 $display("\n2**-487 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2180000000000000;

    #10 $display("\n2**-488 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2170000000000000;

    #10 $display("\n2**-489 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2160000000000000;

    #10 $display("\n2**-490 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2150000000000000;

    #10 $display("\n2**-491 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2140000000000000;

    #10 $display("\n2**-492 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2130000000000000;

    #10 $display("\n2**-493 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2120000000000000;

    #10 $display("\n2**-494 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2110000000000000;

    #10 $display("\n2**-495 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2100000000000000;

    #10 $display("\n2**-496 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h20F0000000000000;

    #10 $display("\n2**-497 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h20E0000000000000;

    #10 $display("\n2**-498 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h20D0000000000000;

    #10 $display("\n2**-499 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h20C0000000000000;

    #10 $display("\n2**-500 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h20B0000000000000;

    #10 $display("\n2**-501 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h20A0000000000000;

    #10 $display("\n2**-502 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2090000000000000;

    #10 $display("\n2**-503 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2080000000000000;

    #10 $display("\n2**-504 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2070000000000000;

    #10 $display("\n2**-505 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2060000000000000;

    #10 $display("\n2**-506 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2050000000000000;

    #10 $display("\n2**-507 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2040000000000000;

    #10 $display("\n2**-508 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2030000000000000;

    #10 $display("\n2**-509 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2020000000000000;

    #10 $display("\n2**-510 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2010000000000000;

    #10 $display("\n2**-511 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h2000000000000000;

    #10 $display("\n2**-512 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1FF0000000000000;

    #10 $display("\n2**-513 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1FE0000000000000;

    #10 $display("\n2**-514 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1FD0000000000000;

    #10 $display("\n2**-515 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1FC0000000000000;

    #10 $display("\n2**-516 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1FB0000000000000;

    #10 $display("\n2**-517 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1FA0000000000000;

    #10 $display("\n2**-518 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1F90000000000000;

    #10 $display("\n2**-519 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1F80000000000000;

    #10 $display("\n2**-520 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1F70000000000000;

    #10 $display("\n2**-521 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1F60000000000000;

    #10 $display("\n2**-522 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1F50000000000000;

    #10 $display("\n2**-523 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1F40000000000000;

    #10 $display("\n2**-524 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1F30000000000000;

    #10 $display("\n2**-525 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1F20000000000000;

    #10 $display("\n2**-526 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1F10000000000000;

    #10 $display("\n2**-527 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1F00000000000000;

    #10 $display("\n2**-528 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1EF0000000000000;

    #10 $display("\n2**-529 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1EE0000000000000;

    #10 $display("\n2**-530 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1ED0000000000000;

    #10 $display("\n2**-531 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1EC0000000000000;

    #10 $display("\n2**-532 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1EB0000000000000;

    #10 $display("\n2**-533 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1EA0000000000000;

    #10 $display("\n2**-534 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1E90000000000000;

    #10 $display("\n2**-535 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1E80000000000000;

    #10 $display("\n2**-536 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1E70000000000000;

    #10 $display("\n2**-537 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1E60000000000000;

    #10 $display("\n2**-538 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1E50000000000000;

    #10 $display("\n2**-539 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1E40000000000000;

    #10 $display("\n2**-540 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1E30000000000000;

    #10 $display("\n2**-541 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1E20000000000000;

    #10 $display("\n2**-542 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1E10000000000000;

    #10 $display("\n2**-543 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1E00000000000000;

    #10 $display("\n2**-544 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1DF0000000000000;

    #10 $display("\n2**-545 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1DE0000000000000;

    #10 $display("\n2**-546 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1DD0000000000000;

    #10 $display("\n2**-547 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1DC0000000000000;

    #10 $display("\n2**-548 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1DB0000000000000;

    #10 $display("\n2**-549 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1DA0000000000000;

    #10 $display("\n2**-550 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1D90000000000000;

    #10 $display("\n2**-551 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1D80000000000000;

    #10 $display("\n2**-552 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1D70000000000000;

    #10 $display("\n2**-553 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1D60000000000000;

    #10 $display("\n2**-554 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1D50000000000000;

    #10 $display("\n2**-555 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1D40000000000000;

    #10 $display("\n2**-556 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1D30000000000000;

    #10 $display("\n2**-557 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1D20000000000000;

    #10 $display("\n2**-558 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1D10000000000000;

    #10 $display("\n2**-559 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1D00000000000000;

    #10 $display("\n2**-560 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1CF0000000000000;

    #10 $display("\n2**-561 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1CE0000000000000;

    #10 $display("\n2**-562 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1CD0000000000000;

    #10 $display("\n2**-563 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1CC0000000000000;

    #10 $display("\n2**-564 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1CB0000000000000;

    #10 $display("\n2**-565 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1CA0000000000000;

    #10 $display("\n2**-566 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1C90000000000000;

    #10 $display("\n2**-567 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1C80000000000000;

    #10 $display("\n2**-568 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1C70000000000000;

    #10 $display("\n2**-569 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1C60000000000000;

    #10 $display("\n2**-570 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1C50000000000000;

    #10 $display("\n2**-571 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1C40000000000000;

    #10 $display("\n2**-572 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1C30000000000000;

    #10 $display("\n2**-573 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1C20000000000000;

    #10 $display("\n2**-574 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1C10000000000000;

    #10 $display("\n2**-575 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1C00000000000000;

    #10 $display("\n2**-576 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1BF0000000000000;

    #10 $display("\n2**-577 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1BE0000000000000;

    #10 $display("\n2**-578 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1BD0000000000000;

    #10 $display("\n2**-579 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1BC0000000000000;

    #10 $display("\n2**-580 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1BB0000000000000;

    #10 $display("\n2**-581 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1BA0000000000000;

    #10 $display("\n2**-582 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1B90000000000000;

    #10 $display("\n2**-583 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1B80000000000000;

    #10 $display("\n2**-584 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1B70000000000000;

    #10 $display("\n2**-585 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1B60000000000000;

    #10 $display("\n2**-586 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1B50000000000000;

    #10 $display("\n2**-587 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1B40000000000000;

    #10 $display("\n2**-588 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1B30000000000000;

    #10 $display("\n2**-589 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1B20000000000000;

    #10 $display("\n2**-590 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1B10000000000000;

    #10 $display("\n2**-591 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1B00000000000000;

    #10 $display("\n2**-592 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1AF0000000000000;

    #10 $display("\n2**-593 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1AE0000000000000;

    #10 $display("\n2**-594 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1AD0000000000000;

    #10 $display("\n2**-595 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1AC0000000000000;

    #10 $display("\n2**-596 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1AB0000000000000;

    #10 $display("\n2**-597 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1AA0000000000000;

    #10 $display("\n2**-598 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1A90000000000000;

    #10 $display("\n2**-599 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1A80000000000000;

    #10 $display("\n2**-600 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1A70000000000000;

    #10 $display("\n2**-601 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1A60000000000000;

    #10 $display("\n2**-602 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1A50000000000000;

    #10 $display("\n2**-603 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1A40000000000000;

    #10 $display("\n2**-604 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1A30000000000000;

    #10 $display("\n2**-605 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1A20000000000000;

    #10 $display("\n2**-606 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1A10000000000000;

    #10 $display("\n2**-607 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1A00000000000000;

    #10 $display("\n2**-608 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h19F0000000000000;

    #10 $display("\n2**-609 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h19E0000000000000;

    #10 $display("\n2**-610 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h19D0000000000000;

    #10 $display("\n2**-611 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h19C0000000000000;

    #10 $display("\n2**-612 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h19B0000000000000;

    #10 $display("\n2**-613 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h19A0000000000000;

    #10 $display("\n2**-614 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1990000000000000;

    #10 $display("\n2**-615 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1980000000000000;

    #10 $display("\n2**-616 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1970000000000000;

    #10 $display("\n2**-617 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1960000000000000;

    #10 $display("\n2**-618 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1950000000000000;

    #10 $display("\n2**-619 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1940000000000000;

    #10 $display("\n2**-620 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1930000000000000;

    #10 $display("\n2**-621 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1920000000000000;

    #10 $display("\n2**-622 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1910000000000000;

    #10 $display("\n2**-623 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1900000000000000;

    #10 $display("\n2**-624 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h18F0000000000000;

    #10 $display("\n2**-625 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h18E0000000000000;

    #10 $display("\n2**-626 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h18D0000000000000;

    #10 $display("\n2**-627 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h18C0000000000000;

    #10 $display("\n2**-628 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h18B0000000000000;

    #10 $display("\n2**-629 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h18A0000000000000;

    #10 $display("\n2**-630 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1890000000000000;

    #10 $display("\n2**-631 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1880000000000000;

    #10 $display("\n2**-632 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1870000000000000;

    #10 $display("\n2**-633 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1860000000000000;

    #10 $display("\n2**-634 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1850000000000000;

    #10 $display("\n2**-635 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1840000000000000;

    #10 $display("\n2**-636 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1830000000000000;

    #10 $display("\n2**-637 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1820000000000000;

    #10 $display("\n2**-638 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1810000000000000;

    #10 $display("\n2**-639 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1800000000000000;

    #10 $display("\n2**-640 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h17F0000000000000;

    #10 $display("\n2**-641 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h17E0000000000000;

    #10 $display("\n2**-642 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h17D0000000000000;

    #10 $display("\n2**-643 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h17C0000000000000;

    #10 $display("\n2**-644 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h17B0000000000000;

    #10 $display("\n2**-645 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h17A0000000000000;

    #10 $display("\n2**-646 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1790000000000000;

    #10 $display("\n2**-647 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1780000000000000;

    #10 $display("\n2**-648 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1770000000000000;

    #10 $display("\n2**-649 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1760000000000000;

    #10 $display("\n2**-650 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1750000000000000;

    #10 $display("\n2**-651 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1740000000000000;

    #10 $display("\n2**-652 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1730000000000000;

    #10 $display("\n2**-653 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1720000000000000;

    #10 $display("\n2**-654 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1710000000000000;

    #10 $display("\n2**-655 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1700000000000000;

    #10 $display("\n2**-656 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h16F0000000000000;

    #10 $display("\n2**-657 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h16E0000000000000;

    #10 $display("\n2**-658 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h16D0000000000000;

    #10 $display("\n2**-659 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h16C0000000000000;

    #10 $display("\n2**-660 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h16B0000000000000;

    #10 $display("\n2**-661 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h16A0000000000000;

    #10 $display("\n2**-662 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1690000000000000;

    #10 $display("\n2**-663 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1680000000000000;

    #10 $display("\n2**-664 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1670000000000000;

    #10 $display("\n2**-665 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1660000000000000;

    #10 $display("\n2**-666 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1650000000000000;

    #10 $display("\n2**-667 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1640000000000000;

    #10 $display("\n2**-668 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1630000000000000;

    #10 $display("\n2**-669 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1620000000000000;

    #10 $display("\n2**-670 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1610000000000000;

    #10 $display("\n2**-671 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1600000000000000;

    #10 $display("\n2**-672 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h15F0000000000000;

    #10 $display("\n2**-673 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h15E0000000000000;

    #10 $display("\n2**-674 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h15D0000000000000;

    #10 $display("\n2**-675 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h15C0000000000000;

    #10 $display("\n2**-676 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h15B0000000000000;

    #10 $display("\n2**-677 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h15A0000000000000;

    #10 $display("\n2**-678 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1590000000000000;

    #10 $display("\n2**-679 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1580000000000000;

    #10 $display("\n2**-680 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1570000000000000;

    #10 $display("\n2**-681 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1560000000000000;

    #10 $display("\n2**-682 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1550000000000000;

    #10 $display("\n2**-683 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1540000000000000;

    #10 $display("\n2**-684 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1530000000000000;

    #10 $display("\n2**-685 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1520000000000000;

    #10 $display("\n2**-686 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1510000000000000;

    #10 $display("\n2**-687 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1500000000000000;

    #10 $display("\n2**-688 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h14F0000000000000;

    #10 $display("\n2**-689 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h14E0000000000000;

    #10 $display("\n2**-690 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h14D0000000000000;

    #10 $display("\n2**-691 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h14C0000000000000;

    #10 $display("\n2**-692 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h14B0000000000000;

    #10 $display("\n2**-693 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h14A0000000000000;

    #10 $display("\n2**-694 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1490000000000000;

    #10 $display("\n2**-695 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1480000000000000;

    #10 $display("\n2**-696 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1470000000000000;

    #10 $display("\n2**-697 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1460000000000000;

    #10 $display("\n2**-698 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1450000000000000;

    #10 $display("\n2**-699 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1440000000000000;

    #10 $display("\n2**-700 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1430000000000000;

    #10 $display("\n2**-701 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1420000000000000;

    #10 $display("\n2**-702 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1410000000000000;

    #10 $display("\n2**-703 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1400000000000000;

    #10 $display("\n2**-704 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h13F0000000000000;

    #10 $display("\n2**-705 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h13E0000000000000;

    #10 $display("\n2**-706 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h13D0000000000000;

    #10 $display("\n2**-707 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h13C0000000000000;

    #10 $display("\n2**-708 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h13B0000000000000;

    #10 $display("\n2**-709 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h13A0000000000000;

    #10 $display("\n2**-710 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1390000000000000;

    #10 $display("\n2**-711 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1380000000000000;

    #10 $display("\n2**-712 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1370000000000000;

    #10 $display("\n2**-713 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1360000000000000;

    #10 $display("\n2**-714 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1350000000000000;

    #10 $display("\n2**-715 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1340000000000000;

    #10 $display("\n2**-716 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1330000000000000;

    #10 $display("\n2**-717 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1320000000000000;

    #10 $display("\n2**-718 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1310000000000000;

    #10 $display("\n2**-719 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1300000000000000;

    #10 $display("\n2**-720 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h12F0000000000000;

    #10 $display("\n2**-721 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h12E0000000000000;

    #10 $display("\n2**-722 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h12D0000000000000;

    #10 $display("\n2**-723 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h12C0000000000000;

    #10 $display("\n2**-724 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h12B0000000000000;

    #10 $display("\n2**-725 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h12A0000000000000;

    #10 $display("\n2**-726 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1290000000000000;

    #10 $display("\n2**-727 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1280000000000000;

    #10 $display("\n2**-728 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1270000000000000;

    #10 $display("\n2**-729 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1260000000000000;

    #10 $display("\n2**-730 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1250000000000000;

    #10 $display("\n2**-731 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1240000000000000;

    #10 $display("\n2**-732 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1230000000000000;

    #10 $display("\n2**-733 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1220000000000000;

    #10 $display("\n2**-734 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1210000000000000;

    #10 $display("\n2**-735 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1200000000000000;

    #10 $display("\n2**-736 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h11F0000000000000;

    #10 $display("\n2**-737 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h11E0000000000000;

    #10 $display("\n2**-738 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h11D0000000000000;

    #10 $display("\n2**-739 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h11C0000000000000;

    #10 $display("\n2**-740 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h11B0000000000000;

    #10 $display("\n2**-741 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h11A0000000000000;

    #10 $display("\n2**-742 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1190000000000000;

    #10 $display("\n2**-743 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1180000000000000;

    #10 $display("\n2**-744 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1170000000000000;

    #10 $display("\n2**-745 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1160000000000000;

    #10 $display("\n2**-746 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1150000000000000;

    #10 $display("\n2**-747 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1140000000000000;

    #10 $display("\n2**-748 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1130000000000000;

    #10 $display("\n2**-749 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1120000000000000;

    #10 $display("\n2**-750 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1110000000000000;

    #10 $display("\n2**-751 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1100000000000000;

    #10 $display("\n2**-752 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h10F0000000000000;

    #10 $display("\n2**-753 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h10E0000000000000;

    #10 $display("\n2**-754 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h10D0000000000000;

    #10 $display("\n2**-755 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h10C0000000000000;

    #10 $display("\n2**-756 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h10B0000000000000;

    #10 $display("\n2**-757 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h10A0000000000000;

    #10 $display("\n2**-758 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1090000000000000;

    #10 $display("\n2**-759 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1080000000000000;

    #10 $display("\n2**-760 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1070000000000000;

    #10 $display("\n2**-761 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1060000000000000;

    #10 $display("\n2**-762 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1050000000000000;

    #10 $display("\n2**-763 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1040000000000000;

    #10 $display("\n2**-764 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1030000000000000;

    #10 $display("\n2**-765 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1020000000000000;

    #10 $display("\n2**-766 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1010000000000000;

    #10 $display("\n2**-767 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h1000000000000000;

    #10 $display("\n2**-768 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0FF0000000000000;

    #10 $display("\n2**-769 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0FE0000000000000;

    #10 $display("\n2**-770 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0FD0000000000000;

    #10 $display("\n2**-771 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0FC0000000000000;

    #10 $display("\n2**-772 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0FB0000000000000;

    #10 $display("\n2**-773 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0FA0000000000000;

    #10 $display("\n2**-774 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0F90000000000000;

    #10 $display("\n2**-775 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0F80000000000000;

    #10 $display("\n2**-776 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0F70000000000000;

    #10 $display("\n2**-777 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0F60000000000000;

    #10 $display("\n2**-778 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0F50000000000000;

    #10 $display("\n2**-779 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0F40000000000000;

    #10 $display("\n2**-780 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0F30000000000000;

    #10 $display("\n2**-781 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0F20000000000000;

    #10 $display("\n2**-782 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0F10000000000000;

    #10 $display("\n2**-783 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0F00000000000000;

    #10 $display("\n2**-784 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0EF0000000000000;

    #10 $display("\n2**-785 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0EE0000000000000;

    #10 $display("\n2**-786 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0ED0000000000000;

    #10 $display("\n2**-787 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0EC0000000000000;

    #10 $display("\n2**-788 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0EB0000000000000;

    #10 $display("\n2**-789 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0EA0000000000000;

    #10 $display("\n2**-790 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0E90000000000000;

    #10 $display("\n2**-791 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0E80000000000000;

    #10 $display("\n2**-792 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0E70000000000000;

    #10 $display("\n2**-793 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0E60000000000000;

    #10 $display("\n2**-794 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0E50000000000000;

    #10 $display("\n2**-795 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0E40000000000000;

    #10 $display("\n2**-796 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0E30000000000000;

    #10 $display("\n2**-797 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0E20000000000000;

    #10 $display("\n2**-798 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0E10000000000000;

    #10 $display("\n2**-799 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0E00000000000000;

    #10 $display("\n2**-800 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0DF0000000000000;

    #10 $display("\n2**-801 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0DE0000000000000;

    #10 $display("\n2**-802 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0DD0000000000000;

    #10 $display("\n2**-803 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0DC0000000000000;

    #10 $display("\n2**-804 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0DB0000000000000;

    #10 $display("\n2**-805 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0DA0000000000000;

    #10 $display("\n2**-806 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0D90000000000000;

    #10 $display("\n2**-807 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0D80000000000000;

    #10 $display("\n2**-808 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0D70000000000000;

    #10 $display("\n2**-809 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0D60000000000000;

    #10 $display("\n2**-810 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0D50000000000000;

    #10 $display("\n2**-811 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0D40000000000000;

    #10 $display("\n2**-812 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0D30000000000000;

    #10 $display("\n2**-813 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0D20000000000000;

    #10 $display("\n2**-814 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0D10000000000000;

    #10 $display("\n2**-815 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0D00000000000000;

    #10 $display("\n2**-816 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0CF0000000000000;

    #10 $display("\n2**-817 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0CE0000000000000;

    #10 $display("\n2**-818 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0CD0000000000000;

    #10 $display("\n2**-819 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0CC0000000000000;

    #10 $display("\n2**-820 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0CB0000000000000;

    #10 $display("\n2**-821 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0CA0000000000000;

    #10 $display("\n2**-822 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0C90000000000000;

    #10 $display("\n2**-823 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0C80000000000000;

    #10 $display("\n2**-824 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0C70000000000000;

    #10 $display("\n2**-825 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0C60000000000000;

    #10 $display("\n2**-826 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0C50000000000000;

    #10 $display("\n2**-827 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0C40000000000000;

    #10 $display("\n2**-828 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0C30000000000000;

    #10 $display("\n2**-829 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0C20000000000000;

    #10 $display("\n2**-830 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0C10000000000000;

    #10 $display("\n2**-831 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0C00000000000000;

    #10 $display("\n2**-832 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0BF0000000000000;

    #10 $display("\n2**-833 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0BE0000000000000;

    #10 $display("\n2**-834 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0BD0000000000000;

    #10 $display("\n2**-835 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0BC0000000000000;

    #10 $display("\n2**-836 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0BB0000000000000;

    #10 $display("\n2**-837 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0BA0000000000000;

    #10 $display("\n2**-838 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0B90000000000000;

    #10 $display("\n2**-839 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0B80000000000000;

    #10 $display("\n2**-840 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0B70000000000000;

    #10 $display("\n2**-841 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0B60000000000000;

    #10 $display("\n2**-842 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0B50000000000000;

    #10 $display("\n2**-843 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0B40000000000000;

    #10 $display("\n2**-844 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0B30000000000000;

    #10 $display("\n2**-845 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0B20000000000000;

    #10 $display("\n2**-846 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0B10000000000000;

    #10 $display("\n2**-847 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0B00000000000000;

    #10 $display("\n2**-848 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0AF0000000000000;

    #10 $display("\n2**-849 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0AE0000000000000;

    #10 $display("\n2**-850 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0AD0000000000000;

    #10 $display("\n2**-851 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0AC0000000000000;

    #10 $display("\n2**-852 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0AB0000000000000;

    #10 $display("\n2**-853 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0AA0000000000000;

    #10 $display("\n2**-854 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0A90000000000000;

    #10 $display("\n2**-855 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0A80000000000000;

    #10 $display("\n2**-856 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0A70000000000000;

    #10 $display("\n2**-857 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0A60000000000000;

    #10 $display("\n2**-858 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0A50000000000000;

    #10 $display("\n2**-859 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0A40000000000000;

    #10 $display("\n2**-860 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0A30000000000000;

    #10 $display("\n2**-861 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0A20000000000000;

    #10 $display("\n2**-862 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0A10000000000000;

    #10 $display("\n2**-863 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0A00000000000000;

    #10 $display("\n2**-864 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h09F0000000000000;

    #10 $display("\n2**-865 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h09E0000000000000;

    #10 $display("\n2**-866 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h09D0000000000000;

    #10 $display("\n2**-867 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h09C0000000000000;

    #10 $display("\n2**-868 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h09B0000000000000;

    #10 $display("\n2**-869 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h09A0000000000000;

    #10 $display("\n2**-870 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0990000000000000;

    #10 $display("\n2**-871 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0980000000000000;

    #10 $display("\n2**-872 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0970000000000000;

    #10 $display("\n2**-873 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0960000000000000;

    #10 $display("\n2**-874 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0950000000000000;

    #10 $display("\n2**-875 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0940000000000000;

    #10 $display("\n2**-876 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0930000000000000;

    #10 $display("\n2**-877 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0920000000000000;

    #10 $display("\n2**-878 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0910000000000000;

    #10 $display("\n2**-879 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0900000000000000;

    #10 $display("\n2**-880 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h08F0000000000000;

    #10 $display("\n2**-881 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h08E0000000000000;

    #10 $display("\n2**-882 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h08D0000000000000;

    #10 $display("\n2**-883 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h08C0000000000000;

    #10 $display("\n2**-884 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h08B0000000000000;

    #10 $display("\n2**-885 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h08A0000000000000;

    #10 $display("\n2**-886 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0890000000000000;

    #10 $display("\n2**-887 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0880000000000000;

    #10 $display("\n2**-888 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0870000000000000;

    #10 $display("\n2**-889 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0860000000000000;

    #10 $display("\n2**-890 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0850000000000000;

    #10 $display("\n2**-891 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0840000000000000;

    #10 $display("\n2**-892 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0830000000000000;

    #10 $display("\n2**-893 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0820000000000000;

    #10 $display("\n2**-894 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0810000000000000;

    #10 $display("\n2**-895 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0800000000000000;

    #10 $display("\n2**-896 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h07F0000000000000;

    #10 $display("\n2**-897 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h07E0000000000000;

    #10 $display("\n2**-898 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h07D0000000000000;

    #10 $display("\n2**-899 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h07C0000000000000;

    #10 $display("\n2**-900 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h07B0000000000000;

    #10 $display("\n2**-901 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h07A0000000000000;

    #10 $display("\n2**-902 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0790000000000000;

    #10 $display("\n2**-903 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0780000000000000;

    #10 $display("\n2**-904 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0770000000000000;

    #10 $display("\n2**-905 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0760000000000000;

    #10 $display("\n2**-906 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0750000000000000;

    #10 $display("\n2**-907 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0740000000000000;

    #10 $display("\n2**-908 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0730000000000000;

    #10 $display("\n2**-909 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0720000000000000;

    #10 $display("\n2**-910 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0710000000000000;

    #10 $display("\n2**-911 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0700000000000000;

    #10 $display("\n2**-912 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h06F0000000000000;

    #10 $display("\n2**-913 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h06E0000000000000;

    #10 $display("\n2**-914 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h06D0000000000000;

    #10 $display("\n2**-915 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h06C0000000000000;

    #10 $display("\n2**-916 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h06B0000000000000;

    #10 $display("\n2**-917 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h06A0000000000000;

    #10 $display("\n2**-918 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0690000000000000;

    #10 $display("\n2**-919 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0680000000000000;

    #10 $display("\n2**-920 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0670000000000000;

    #10 $display("\n2**-921 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0660000000000000;

    #10 $display("\n2**-922 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0650000000000000;

    #10 $display("\n2**-923 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0640000000000000;

    #10 $display("\n2**-924 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0630000000000000;

    #10 $display("\n2**-925 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0620000000000000;

    #10 $display("\n2**-926 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0610000000000000;

    #10 $display("\n2**-927 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0600000000000000;

    #10 $display("\n2**-928 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h05F0000000000000;

    #10 $display("\n2**-929 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h05E0000000000000;

    #10 $display("\n2**-930 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h05D0000000000000;

    #10 $display("\n2**-931 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h05C0000000000000;

    #10 $display("\n2**-932 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h05B0000000000000;

    #10 $display("\n2**-933 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h05A0000000000000;

    #10 $display("\n2**-934 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0590000000000000;

    #10 $display("\n2**-935 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0580000000000000;

    #10 $display("\n2**-936 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0570000000000000;

    #10 $display("\n2**-937 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0560000000000000;

    #10 $display("\n2**-938 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0550000000000000;

    #10 $display("\n2**-939 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0540000000000000;

    #10 $display("\n2**-940 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0530000000000000;

    #10 $display("\n2**-941 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0520000000000000;

    #10 $display("\n2**-942 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0510000000000000;

    #10 $display("\n2**-943 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0500000000000000;

    #10 $display("\n2**-944 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h04F0000000000000;

    #10 $display("\n2**-945 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h04E0000000000000;

    #10 $display("\n2**-946 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h04D0000000000000;

    #10 $display("\n2**-947 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h04C0000000000000;

    #10 $display("\n2**-948 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h04B0000000000000;

    #10 $display("\n2**-949 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h04A0000000000000;

    #10 $display("\n2**-950 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0490000000000000;

    #10 $display("\n2**-951 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0480000000000000;

    #10 $display("\n2**-952 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0470000000000000;

    #10 $display("\n2**-953 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0460000000000000;

    #10 $display("\n2**-954 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0450000000000000;

    #10 $display("\n2**-955 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0440000000000000;

    #10 $display("\n2**-956 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0430000000000000;

    #10 $display("\n2**-957 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0420000000000000;

    #10 $display("\n2**-958 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0410000000000000;

    #10 $display("\n2**-959 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0400000000000000;

    #10 $display("\n2**-960 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h03F0000000000000;

    #10 $display("\n2**-961 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h03E0000000000000;

    #10 $display("\n2**-962 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h03D0000000000000;

    #10 $display("\n2**-963 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h03C0000000000000;

    #10 $display("\n2**-964 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h03B0000000000000;

    #10 $display("\n2**-965 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h03A0000000000000;

    #10 $display("\n2**-966 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0390000000000000;

    #10 $display("\n2**-967 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0380000000000000;

    #10 $display("\n2**-968 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0370000000000000;

    #10 $display("\n2**-969 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0360000000000000;

    #10 $display("\n2**-970 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0350000000000000;

    #10 $display("\n2**-971 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0340000000000000;

    #10 $display("\n2**-972 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0330000000000000;

    #10 $display("\n2**-973 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0320000000000000;

    #10 $display("\n2**-974 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0310000000000000;

    #10 $display("\n2**-975 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0300000000000000;

    #10 $display("\n2**-976 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h02F0000000000000;

    #10 $display("\n2**-977 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h02E0000000000000;

    #10 $display("\n2**-978 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h02D0000000000000;

    #10 $display("\n2**-979 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h02C0000000000000;

    #10 $display("\n2**-980 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h02B0000000000000;

    #10 $display("\n2**-981 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h02A0000000000000;

    #10 $display("\n2**-982 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0290000000000000;

    #10 $display("\n2**-983 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0280000000000000;

    #10 $display("\n2**-984 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0270000000000000;

    #10 $display("\n2**-985 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0260000000000000;

    #10 $display("\n2**-986 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0250000000000000;

    #10 $display("\n2**-987 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0240000000000000;

    #10 $display("\n2**-988 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0230000000000000;

    #10 $display("\n2**-989 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0220000000000000;

    #10 $display("\n2**-990 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0210000000000000;

    #10 $display("\n2**-991 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0200000000000000;

    #10 $display("\n2**-992 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h01F0000000000000;

    #10 $display("\n2**-993 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h01E0000000000000;

    #10 $display("\n2**-994 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h01D0000000000000;

    #10 $display("\n2**-995 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h01C0000000000000;

    #10 $display("\n2**-996 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h01B0000000000000;

    #10 $display("\n2**-997 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h01A0000000000000;

    #10 $display("\n2**-998 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0190000000000000;

    #10 $display("\n2**-999 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0180000000000000;

    #10 $display("\n2**-1000 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0170000000000000;

    #10 $display("\n2**-1001 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0160000000000000;

    #10 $display("\n2**-1002 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0150000000000000;

    #10 $display("\n2**-1003 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0140000000000000;

    #10 $display("\n2**-1004 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0130000000000000;

    #10 $display("\n2**-1005 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0120000000000000;

    #10 $display("\n2**-1006 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0110000000000000;

    #10 $display("\n2**-1007 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0100000000000000;

    #10 $display("\n2**-1008 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h00F0000000000000;

    #10 $display("\n2**-1009 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h00E0000000000000;

    #10 $display("\n2**-1010 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h00D0000000000000;

    #10 $display("\n2**-1011 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h00C0000000000000;

    #10 $display("\n2**-1012 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h00B0000000000000;

    #10 $display("\n2**-1013 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h00A0000000000000;

    #10 $display("\n2**-1014 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0090000000000000;

    #10 $display("\n2**-1015 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0080000000000000;

    #10 $display("\n2**-1016 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0070000000000000;

    #10 $display("\n2**-1017 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0060000000000000;

    #10 $display("\n2**-1018 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0050000000000000;

    #10 $display("\n2**-1019 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0040000000000000;

    #10 $display("\n2**-1020 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0030000000000000;

    #10 $display("\n2**-1021 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0020000000000000;

    #10 $display("\n2**-1022 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0010000000000000;

    #10 $display("\n2**-1023 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0008000000000000;

    #10 $display("\n2**-1024 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0004000000000000;

    #10 $display("\n2**-1025 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0002000000000000;

    #10 $display("\n2**-1026 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0001000000000000;

    #10 $display("\n2**-1027 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000800000000000;

    #10 $display("\n2**-1028 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000400000000000;

    #10 $display("\n2**-1029 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000200000000000;

    #10 $display("\n2**-1030 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000100000000000;

    #10 $display("\n2**-1031 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000080000000000;

    #10 $display("\n2**-1032 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000040000000000;

    #10 $display("\n2**-1033 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000020000000000;

    #10 $display("\n2**-1034 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000010000000000;

    #10 $display("\n2**-1035 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000008000000000;

    #10 $display("\n2**-1036 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000004000000000;

    #10 $display("\n2**-1037 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000002000000000;

    #10 $display("\n2**-1038 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000001000000000;

    #10 $display("\n2**-1039 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000800000000;

    #10 $display("\n2**-1040 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000400000000;

    #10 $display("\n2**-1041 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000200000000;

    #10 $display("\n2**-1042 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000100000000;

    #10 $display("\n2**-1043 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000080000000;

    #10 $display("\n2**-1044 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000040000000;

    #10 $display("\n2**-1045 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000020000000;

    #10 $display("\n2**-1046 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000010000000;

    #10 $display("\n2**-1047 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000008000000;

    #10 $display("\n2**-1048 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000004000000;

    #10 $display("\n2**-1049 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000002000000;

    #10 $display("\n2**-1050 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000001000000;

    #10 $display("\n2**-1051 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000800000;

    #10 $display("\n2**-1052 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000400000;

    #10 $display("\n2**-1053 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000200000;

    #10 $display("\n2**-1054 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000100000;

    #10 $display("\n2**-1055 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000080000;

    #10 $display("\n2**-1056 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000040000;

    #10 $display("\n2**-1057 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000020000;

    #10 $display("\n2**-1058 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000010000;

    #10 $display("\n2**-1059 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000008000;

    #10 $display("\n2**-1060 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000004000;

    #10 $display("\n2**-1061 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000002000;

    #10 $display("\n2**-1062 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000001000;

    #10 $display("\n2**-1063 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000000800;

    #10 $display("\n2**-1064 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000000400;

    #10 $display("\n2**-1065 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000000200;

    #10 $display("\n2**-1066 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000000100;

    #10 $display("\n2**-1067 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000000080;

    #10 $display("\n2**-1068 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000000040;

    #10 $display("\n2**-1069 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000000020;

    #10 $display("\n2**-1070 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000000010;

    #10 $display("\n2**-1071 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000000008;

    #10 $display("\n2**-1072 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000000004;

    #10 $display("\n2**-1073 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000000002;

    #10 $display("\n2**-1074 * 1:");
    #10 assign b = 64'h3FF0000000000000; assign a = 64'h0000000000000001;

    #10 $display("\n2**0 * 2**1023:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h7FE0000000000000;
    #10 assign a = 64'h3FFFFFFFFFFFFFFF; assign b = 64'h7FEFFFFFFFFFFFFF;

    #10 $display("\n2**1 * 2**1022:");
    #10 assign a = 64'h4000000000000000; assign b = 64'h7FD0000000000000;
    #10 assign a = 64'h400FFFFFFFFFFFFF; assign b = 64'h7FDFFFFFFFFFFFFF;

    #10 $display("\n2**2 * 2**1021:");
    #10 assign a = 64'h4010000000000000; assign b = 64'h7FC0000000000000;
    #10 assign a = 64'h401FFFFFFFFFFFFF; assign b = 64'h7FCFFFFFFFFFFFFF;

    #10 $display("\n2**3 * 2**1020:");
    #10 assign a = 64'h4020000000000000; assign b = 64'h7FB0000000000000;
    #10 assign a = 64'h402FFFFFFFFFFFFF; assign b = 64'h7FBFFFFFFFFFFFFF;

    #10 $display("\n2**4 * 2**1019:");
    #10 assign a = 64'h4030000000000000; assign b = 64'h7FA0000000000000;
    #10 assign a = 64'h403FFFFFFFFFFFFF; assign b = 64'h7FAFFFFFFFFFFFFF;

    #10 $display("\n2**5 * 2**1018:");
    #10 assign a = 64'h4040000000000000; assign b = 64'h7F90000000000000;
    #10 assign a = 64'h404FFFFFFFFFFFFF; assign b = 64'h7F9FFFFFFFFFFFFF;

    #10 $display("\n2**6 * 2**1017:");
    #10 assign a = 64'h4050000000000000; assign b = 64'h7F80000000000000;
    #10 assign a = 64'h405FFFFFFFFFFFFF; assign b = 64'h7F8FFFFFFFFFFFFF;

    #10 $display("\n2**7 * 2**1016:");
    #10 assign a = 64'h4060000000000000; assign b = 64'h7F70000000000000;
    #10 assign a = 64'h406FFFFFFFFFFFFF; assign b = 64'h7F7FFFFFFFFFFFFF;

    #10 $display("\n2**8 * 2**1015:");
    #10 assign a = 64'h4070000000000000; assign b = 64'h7F60000000000000;
    #10 assign a = 64'h407FFFFFFFFFFFFF; assign b = 64'h7F6FFFFFFFFFFFFF;

    #10 $display("\n2**9 * 2**1014:");
    #10 assign a = 64'h4080000000000000; assign b = 64'h7F50000000000000;
    #10 assign a = 64'h408FFFFFFFFFFFFF; assign b = 64'h7F5FFFFFFFFFFFFF;

    #10 $display("\n2**10 * 2**1013:");
    #10 assign a = 64'h4090000000000000; assign b = 64'h7F40000000000000;
    #10 assign a = 64'h409FFFFFFFFFFFFF; assign b = 64'h7F4FFFFFFFFFFFFF;

    #10 $display("\n2**11 * 2**1012:");
    #10 assign a = 64'h40A0000000000000; assign b = 64'h7F30000000000000;
    #10 assign a = 64'h40AFFFFFFFFFFFFF; assign b = 64'h7F3FFFFFFFFFFFFF;

    #10 $display("\n2**12 * 2**1011:");
    #10 assign a = 64'h40B0000000000000; assign b = 64'h7F20000000000000;
    #10 assign a = 64'h40BFFFFFFFFFFFFF; assign b = 64'h7F2FFFFFFFFFFFFF;

    #10 $display("\n2**13 * 2**1010:");
    #10 assign a = 64'h40C0000000000000; assign b = 64'h7F10000000000000;
    #10 assign a = 64'h40CFFFFFFFFFFFFF; assign b = 64'h7F1FFFFFFFFFFFFF;

    #10 $display("\n2**14 * 2**1009:");
    #10 assign a = 64'h40D0000000000000; assign b = 64'h7F00000000000000;
    #10 assign a = 64'h40DFFFFFFFFFFFFF; assign b = 64'h7F0FFFFFFFFFFFFF;

    #10 $display("\n2**15 * 2**1008:");
    #10 assign a = 64'h40E0000000000000; assign b = 64'h7EF0000000000000;
    #10 assign a = 64'h40EFFFFFFFFFFFFF; assign b = 64'h7EFFFFFFFFFFFFFF;

    #10 $display("\n2**16 * 2**1007:");
    #10 assign a = 64'h40F0000000000000; assign b = 64'h7EE0000000000000;
    #10 assign a = 64'h40FFFFFFFFFFFFFF; assign b = 64'h7EEFFFFFFFFFFFFF;

    #10 $display("\n2**17 * 2**1006:");
    #10 assign a = 64'h4100000000000000; assign b = 64'h7ED0000000000000;
    #10 assign a = 64'h410FFFFFFFFFFFFF; assign b = 64'h7EDFFFFFFFFFFFFF;

    #10 $display("\n2**18 * 2**1005:");
    #10 assign a = 64'h4110000000000000; assign b = 64'h7EC0000000000000;
    #10 assign a = 64'h411FFFFFFFFFFFFF; assign b = 64'h7ECFFFFFFFFFFFFF;

    #10 $display("\n2**19 * 2**1004:");
    #10 assign a = 64'h4120000000000000; assign b = 64'h7EB0000000000000;
    #10 assign a = 64'h412FFFFFFFFFFFFF; assign b = 64'h7EBFFFFFFFFFFFFF;

    #10 $display("\n2**20 * 2**1003:");
    #10 assign a = 64'h4130000000000000; assign b = 64'h7EA0000000000000;
    #10 assign a = 64'h413FFFFFFFFFFFFF; assign b = 64'h7EAFFFFFFFFFFFFF;

    #10 $display("\n2**21 * 2**1002:");
    #10 assign a = 64'h4140000000000000; assign b = 64'h7E90000000000000;
    #10 assign a = 64'h414FFFFFFFFFFFFF; assign b = 64'h7E9FFFFFFFFFFFFF;

    #10 $display("\n2**22 * 2**1001:");
    #10 assign a = 64'h4150000000000000; assign b = 64'h7E80000000000000;
    #10 assign a = 64'h415FFFFFFFFFFFFF; assign b = 64'h7E8FFFFFFFFFFFFF;

    #10 $display("\n2**23 * 2**1000:");
    #10 assign a = 64'h4160000000000000; assign b = 64'h7E70000000000000;
    #10 assign a = 64'h416FFFFFFFFFFFFF; assign b = 64'h7E7FFFFFFFFFFFFF;

    #10 $display("\n2**24 * 2**999:");
    #10 assign a = 64'h4170000000000000; assign b = 64'h7E60000000000000;
    #10 assign a = 64'h417FFFFFFFFFFFFF; assign b = 64'h7E6FFFFFFFFFFFFF;

    #10 $display("\n2**25 * 2**998:");
    #10 assign a = 64'h4180000000000000; assign b = 64'h7E50000000000000;
    #10 assign a = 64'h418FFFFFFFFFFFFF; assign b = 64'h7E5FFFFFFFFFFFFF;

    #10 $display("\n2**26 * 2**997:");
    #10 assign a = 64'h4190000000000000; assign b = 64'h7E40000000000000;
    #10 assign a = 64'h419FFFFFFFFFFFFF; assign b = 64'h7E4FFFFFFFFFFFFF;

    #10 $display("\n2**27 * 2**996:");
    #10 assign a = 64'h41A0000000000000; assign b = 64'h7E30000000000000;
    #10 assign a = 64'h41AFFFFFFFFFFFFF; assign b = 64'h7E3FFFFFFFFFFFFF;

    #10 $display("\n2**28 * 2**995:");
    #10 assign a = 64'h41B0000000000000; assign b = 64'h7E20000000000000;
    #10 assign a = 64'h41BFFFFFFFFFFFFF; assign b = 64'h7E2FFFFFFFFFFFFF;

    #10 $display("\n2**29 * 2**994:");
    #10 assign a = 64'h41C0000000000000; assign b = 64'h7E10000000000000;
    #10 assign a = 64'h41CFFFFFFFFFFFFF; assign b = 64'h7E1FFFFFFFFFFFFF;

    #10 $display("\n2**30 * 2**993:");
    #10 assign a = 64'h41D0000000000000; assign b = 64'h7E00000000000000;
    #10 assign a = 64'h41DFFFFFFFFFFFFF; assign b = 64'h7E0FFFFFFFFFFFFF;

    #10 $display("\n2**31 * 2**992:");
    #10 assign a = 64'h41E0000000000000; assign b = 64'h7DF0000000000000;
    #10 assign a = 64'h41EFFFFFFFFFFFFF; assign b = 64'h7DFFFFFFFFFFFFFF;

    #10 $display("\n2**32 * 2**991:");
    #10 assign a = 64'h41F0000000000000; assign b = 64'h7DE0000000000000;
    #10 assign a = 64'h41FFFFFFFFFFFFFF; assign b = 64'h7DEFFFFFFFFFFFFF;

    #10 $display("\n2**33 * 2**990:");
    #10 assign a = 64'h4200000000000000; assign b = 64'h7DD0000000000000;
    #10 assign a = 64'h420FFFFFFFFFFFFF; assign b = 64'h7DDFFFFFFFFFFFFF;

    #10 $display("\n2**34 * 2**989:");
    #10 assign a = 64'h4210000000000000; assign b = 64'h7DC0000000000000;
    #10 assign a = 64'h421FFFFFFFFFFFFF; assign b = 64'h7DCFFFFFFFFFFFFF;

    #10 $display("\n2**35 * 2**988:");
    #10 assign a = 64'h4220000000000000; assign b = 64'h7DB0000000000000;
    #10 assign a = 64'h422FFFFFFFFFFFFF; assign b = 64'h7DBFFFFFFFFFFFFF;

    #10 $display("\n2**36 * 2**987:");
    #10 assign a = 64'h4230000000000000; assign b = 64'h7DA0000000000000;
    #10 assign a = 64'h423FFFFFFFFFFFFF; assign b = 64'h7DAFFFFFFFFFFFFF;

    #10 $display("\n2**37 * 2**986:");
    #10 assign a = 64'h4240000000000000; assign b = 64'h7D90000000000000;
    #10 assign a = 64'h424FFFFFFFFFFFFF; assign b = 64'h7D9FFFFFFFFFFFFF;

    #10 $display("\n2**38 * 2**985:");
    #10 assign a = 64'h4250000000000000; assign b = 64'h7D80000000000000;
    #10 assign a = 64'h425FFFFFFFFFFFFF; assign b = 64'h7D8FFFFFFFFFFFFF;

    #10 $display("\n2**39 * 2**984:");
    #10 assign a = 64'h4260000000000000; assign b = 64'h7D70000000000000;
    #10 assign a = 64'h426FFFFFFFFFFFFF; assign b = 64'h7D7FFFFFFFFFFFFF;

    #10 $display("\n2**40 * 2**983:");
    #10 assign a = 64'h4270000000000000; assign b = 64'h7D60000000000000;
    #10 assign a = 64'h427FFFFFFFFFFFFF; assign b = 64'h7D6FFFFFFFFFFFFF;

    #10 $display("\n2**41 * 2**982:");
    #10 assign a = 64'h4280000000000000; assign b = 64'h7D50000000000000;
    #10 assign a = 64'h428FFFFFFFFFFFFF; assign b = 64'h7D5FFFFFFFFFFFFF;

    #10 $display("\n2**42 * 2**981:");
    #10 assign a = 64'h4290000000000000; assign b = 64'h7D40000000000000;
    #10 assign a = 64'h429FFFFFFFFFFFFF; assign b = 64'h7D4FFFFFFFFFFFFF;

    #10 $display("\n2**43 * 2**980:");
    #10 assign a = 64'h42A0000000000000; assign b = 64'h7D30000000000000;
    #10 assign a = 64'h42AFFFFFFFFFFFFF; assign b = 64'h7D3FFFFFFFFFFFFF;

    #10 $display("\n2**44 * 2**979:");
    #10 assign a = 64'h42B0000000000000; assign b = 64'h7D20000000000000;
    #10 assign a = 64'h42BFFFFFFFFFFFFF; assign b = 64'h7D2FFFFFFFFFFFFF;

    #10 $display("\n2**45 * 2**978:");
    #10 assign a = 64'h42C0000000000000; assign b = 64'h7D10000000000000;
    #10 assign a = 64'h42CFFFFFFFFFFFFF; assign b = 64'h7D1FFFFFFFFFFFFF;

    #10 $display("\n2**46 * 2**977:");
    #10 assign a = 64'h42D0000000000000; assign b = 64'h7D00000000000000;
    #10 assign a = 64'h42DFFFFFFFFFFFFF; assign b = 64'h7D0FFFFFFFFFFFFF;

    #10 $display("\n2**47 * 2**976:");
    #10 assign a = 64'h42E0000000000000; assign b = 64'h7CF0000000000000;
    #10 assign a = 64'h42EFFFFFFFFFFFFF; assign b = 64'h7CFFFFFFFFFFFFFF;

    #10 $display("\n2**48 * 2**975:");
    #10 assign a = 64'h42F0000000000000; assign b = 64'h7CE0000000000000;
    #10 assign a = 64'h42FFFFFFFFFFFFFF; assign b = 64'h7CEFFFFFFFFFFFFF;

    #10 $display("\n2**49 * 2**974:");
    #10 assign a = 64'h4300000000000000; assign b = 64'h7CD0000000000000;
    #10 assign a = 64'h430FFFFFFFFFFFFF; assign b = 64'h7CDFFFFFFFFFFFFF;

    #10 $display("\n2**50 * 2**973:");
    #10 assign a = 64'h4310000000000000; assign b = 64'h7CC0000000000000;
    #10 assign a = 64'h431FFFFFFFFFFFFF; assign b = 64'h7CCFFFFFFFFFFFFF;

    #10 $display("\n2**51 * 2**972:");
    #10 assign a = 64'h4320000000000000; assign b = 64'h7CB0000000000000;
    #10 assign a = 64'h432FFFFFFFFFFFFF; assign b = 64'h7CBFFFFFFFFFFFFF;

    #10 $display("\n2**52 * 2**971:");
    #10 assign a = 64'h4330000000000000; assign b = 64'h7CA0000000000000;
    #10 assign a = 64'h433FFFFFFFFFFFFF; assign b = 64'h7CAFFFFFFFFFFFFF;

    #10 $display("\n2**53 * 2**970:");
    #10 assign a = 64'h4340000000000000; assign b = 64'h7C90000000000000;
    #10 assign a = 64'h434FFFFFFFFFFFFF; assign b = 64'h7C9FFFFFFFFFFFFF;

    #10 $display("\n2**54 * 2**969:");
    #10 assign a = 64'h4350000000000000; assign b = 64'h7C80000000000000;
    #10 assign a = 64'h435FFFFFFFFFFFFF; assign b = 64'h7C8FFFFFFFFFFFFF;

    #10 $display("\n2**55 * 2**968:");
    #10 assign a = 64'h4360000000000000; assign b = 64'h7C70000000000000;
    #10 assign a = 64'h436FFFFFFFFFFFFF; assign b = 64'h7C7FFFFFFFFFFFFF;

    #10 $display("\n2**56 * 2**967:");
    #10 assign a = 64'h4370000000000000; assign b = 64'h7C60000000000000;
    #10 assign a = 64'h437FFFFFFFFFFFFF; assign b = 64'h7C6FFFFFFFFFFFFF;

    #10 $display("\n2**57 * 2**966:");
    #10 assign a = 64'h4380000000000000; assign b = 64'h7C50000000000000;
    #10 assign a = 64'h438FFFFFFFFFFFFF; assign b = 64'h7C5FFFFFFFFFFFFF;

    #10 $display("\n2**58 * 2**965:");
    #10 assign a = 64'h4390000000000000; assign b = 64'h7C40000000000000;
    #10 assign a = 64'h439FFFFFFFFFFFFF; assign b = 64'h7C4FFFFFFFFFFFFF;

    #10 $display("\n2**59 * 2**964:");
    #10 assign a = 64'h43A0000000000000; assign b = 64'h7C30000000000000;
    #10 assign a = 64'h43AFFFFFFFFFFFFF; assign b = 64'h7C3FFFFFFFFFFFFF;

    #10 $display("\n2**60 * 2**963:");
    #10 assign a = 64'h43B0000000000000; assign b = 64'h7C20000000000000;
    #10 assign a = 64'h43BFFFFFFFFFFFFF; assign b = 64'h7C2FFFFFFFFFFFFF;

    #10 $display("\n2**61 * 2**962:");
    #10 assign a = 64'h43C0000000000000; assign b = 64'h7C10000000000000;
    #10 assign a = 64'h43CFFFFFFFFFFFFF; assign b = 64'h7C1FFFFFFFFFFFFF;

    #10 $display("\n2**62 * 2**961:");
    #10 assign a = 64'h43D0000000000000; assign b = 64'h7C00000000000000;
    #10 assign a = 64'h43DFFFFFFFFFFFFF; assign b = 64'h7C0FFFFFFFFFFFFF;

    #10 $display("\n2**63 * 2**960:");
    #10 assign a = 64'h43E0000000000000; assign b = 64'h7BF0000000000000;
    #10 assign a = 64'h43EFFFFFFFFFFFFF; assign b = 64'h7BFFFFFFFFFFFFFF;

    #10 $display("\n2**64 * 2**959:");
    #10 assign a = 64'h43F0000000000000; assign b = 64'h7BE0000000000000;
    #10 assign a = 64'h43FFFFFFFFFFFFFF; assign b = 64'h7BEFFFFFFFFFFFFF;

    #10 $display("\n2**65 * 2**958:");
    #10 assign a = 64'h4400000000000000; assign b = 64'h7BD0000000000000;
    #10 assign a = 64'h440FFFFFFFFFFFFF; assign b = 64'h7BDFFFFFFFFFFFFF;

    #10 $display("\n2**66 * 2**957:");
    #10 assign a = 64'h4410000000000000; assign b = 64'h7BC0000000000000;
    #10 assign a = 64'h441FFFFFFFFFFFFF; assign b = 64'h7BCFFFFFFFFFFFFF;

    #10 $display("\n2**67 * 2**956:");
    #10 assign a = 64'h4420000000000000; assign b = 64'h7BB0000000000000;
    #10 assign a = 64'h442FFFFFFFFFFFFF; assign b = 64'h7BBFFFFFFFFFFFFF;

    #10 $display("\n2**68 * 2**955:");
    #10 assign a = 64'h4430000000000000; assign b = 64'h7BA0000000000000;
    #10 assign a = 64'h443FFFFFFFFFFFFF; assign b = 64'h7BAFFFFFFFFFFFFF;

    #10 $display("\n2**69 * 2**954:");
    #10 assign a = 64'h4440000000000000; assign b = 64'h7B90000000000000;
    #10 assign a = 64'h444FFFFFFFFFFFFF; assign b = 64'h7B9FFFFFFFFFFFFF;

    #10 $display("\n2**70 * 2**953:");
    #10 assign a = 64'h4450000000000000; assign b = 64'h7B80000000000000;
    #10 assign a = 64'h445FFFFFFFFFFFFF; assign b = 64'h7B8FFFFFFFFFFFFF;

    #10 $display("\n2**71 * 2**952:");
    #10 assign a = 64'h4460000000000000; assign b = 64'h7B70000000000000;
    #10 assign a = 64'h446FFFFFFFFFFFFF; assign b = 64'h7B7FFFFFFFFFFFFF;

    #10 $display("\n2**72 * 2**951:");
    #10 assign a = 64'h4470000000000000; assign b = 64'h7B60000000000000;
    #10 assign a = 64'h447FFFFFFFFFFFFF; assign b = 64'h7B6FFFFFFFFFFFFF;

    #10 $display("\n2**73 * 2**950:");
    #10 assign a = 64'h4480000000000000; assign b = 64'h7B50000000000000;
    #10 assign a = 64'h448FFFFFFFFFFFFF; assign b = 64'h7B5FFFFFFFFFFFFF;

    #10 $display("\n2**74 * 2**949:");
    #10 assign a = 64'h4490000000000000; assign b = 64'h7B40000000000000;
    #10 assign a = 64'h449FFFFFFFFFFFFF; assign b = 64'h7B4FFFFFFFFFFFFF;

    #10 $display("\n2**75 * 2**948:");
    #10 assign a = 64'h44A0000000000000; assign b = 64'h7B30000000000000;
    #10 assign a = 64'h44AFFFFFFFFFFFFF; assign b = 64'h7B3FFFFFFFFFFFFF;

    #10 $display("\n2**76 * 2**947:");
    #10 assign a = 64'h44B0000000000000; assign b = 64'h7B20000000000000;
    #10 assign a = 64'h44BFFFFFFFFFFFFF; assign b = 64'h7B2FFFFFFFFFFFFF;

    #10 $display("\n2**77 * 2**946:");
    #10 assign a = 64'h44C0000000000000; assign b = 64'h7B10000000000000;
    #10 assign a = 64'h44CFFFFFFFFFFFFF; assign b = 64'h7B1FFFFFFFFFFFFF;

    #10 $display("\n2**78 * 2**945:");
    #10 assign a = 64'h44D0000000000000; assign b = 64'h7B00000000000000;
    #10 assign a = 64'h44DFFFFFFFFFFFFF; assign b = 64'h7B0FFFFFFFFFFFFF;

    #10 $display("\n2**79 * 2**944:");
    #10 assign a = 64'h44E0000000000000; assign b = 64'h7AF0000000000000;
    #10 assign a = 64'h44EFFFFFFFFFFFFF; assign b = 64'h7AFFFFFFFFFFFFFF;

    #10 $display("\n2**80 * 2**943:");
    #10 assign a = 64'h44F0000000000000; assign b = 64'h7AE0000000000000;
    #10 assign a = 64'h44FFFFFFFFFFFFFF; assign b = 64'h7AEFFFFFFFFFFFFF;

    #10 $display("\n2**81 * 2**942:");
    #10 assign a = 64'h4500000000000000; assign b = 64'h7AD0000000000000;
    #10 assign a = 64'h450FFFFFFFFFFFFF; assign b = 64'h7ADFFFFFFFFFFFFF;

    #10 $display("\n2**82 * 2**941:");
    #10 assign a = 64'h4510000000000000; assign b = 64'h7AC0000000000000;
    #10 assign a = 64'h451FFFFFFFFFFFFF; assign b = 64'h7ACFFFFFFFFFFFFF;

    #10 $display("\n2**83 * 2**940:");
    #10 assign a = 64'h4520000000000000; assign b = 64'h7AB0000000000000;
    #10 assign a = 64'h452FFFFFFFFFFFFF; assign b = 64'h7ABFFFFFFFFFFFFF;

    #10 $display("\n2**84 * 2**939:");
    #10 assign a = 64'h4530000000000000; assign b = 64'h7AA0000000000000;
    #10 assign a = 64'h453FFFFFFFFFFFFF; assign b = 64'h7AAFFFFFFFFFFFFF;

    #10 $display("\n2**85 * 2**938:");
    #10 assign a = 64'h4540000000000000; assign b = 64'h7A90000000000000;
    #10 assign a = 64'h454FFFFFFFFFFFFF; assign b = 64'h7A9FFFFFFFFFFFFF;

    #10 $display("\n2**86 * 2**937:");
    #10 assign a = 64'h4550000000000000; assign b = 64'h7A80000000000000;
    #10 assign a = 64'h455FFFFFFFFFFFFF; assign b = 64'h7A8FFFFFFFFFFFFF;

    #10 $display("\n2**87 * 2**936:");
    #10 assign a = 64'h4560000000000000; assign b = 64'h7A70000000000000;
    #10 assign a = 64'h456FFFFFFFFFFFFF; assign b = 64'h7A7FFFFFFFFFFFFF;

    #10 $display("\n2**88 * 2**935:");
    #10 assign a = 64'h4570000000000000; assign b = 64'h7A60000000000000;
    #10 assign a = 64'h457FFFFFFFFFFFFF; assign b = 64'h7A6FFFFFFFFFFFFF;

    #10 $display("\n2**89 * 2**934:");
    #10 assign a = 64'h4580000000000000; assign b = 64'h7A50000000000000;
    #10 assign a = 64'h458FFFFFFFFFFFFF; assign b = 64'h7A5FFFFFFFFFFFFF;

    #10 $display("\n2**90 * 2**933:");
    #10 assign a = 64'h4590000000000000; assign b = 64'h7A40000000000000;
    #10 assign a = 64'h459FFFFFFFFFFFFF; assign b = 64'h7A4FFFFFFFFFFFFF;

    #10 $display("\n2**91 * 2**932:");
    #10 assign a = 64'h45A0000000000000; assign b = 64'h7A30000000000000;
    #10 assign a = 64'h45AFFFFFFFFFFFFF; assign b = 64'h7A3FFFFFFFFFFFFF;

    #10 $display("\n2**92 * 2**931:");
    #10 assign a = 64'h45B0000000000000; assign b = 64'h7A20000000000000;
    #10 assign a = 64'h45BFFFFFFFFFFFFF; assign b = 64'h7A2FFFFFFFFFFFFF;

    #10 $display("\n2**93 * 2**930:");
    #10 assign a = 64'h45C0000000000000; assign b = 64'h7A10000000000000;
    #10 assign a = 64'h45CFFFFFFFFFFFFF; assign b = 64'h7A1FFFFFFFFFFFFF;

    #10 $display("\n2**94 * 2**929:");
    #10 assign a = 64'h45D0000000000000; assign b = 64'h7A00000000000000;
    #10 assign a = 64'h45DFFFFFFFFFFFFF; assign b = 64'h7A0FFFFFFFFFFFFF;

    #10 $display("\n2**95 * 2**928:");
    #10 assign a = 64'h45E0000000000000; assign b = 64'h79F0000000000000;
    #10 assign a = 64'h45EFFFFFFFFFFFFF; assign b = 64'h79FFFFFFFFFFFFFF;

    #10 $display("\n2**96 * 2**927:");
    #10 assign a = 64'h45F0000000000000; assign b = 64'h79E0000000000000;
    #10 assign a = 64'h45FFFFFFFFFFFFFF; assign b = 64'h79EFFFFFFFFFFFFF;

    #10 $display("\n2**97 * 2**926:");
    #10 assign a = 64'h4600000000000000; assign b = 64'h79D0000000000000;
    #10 assign a = 64'h460FFFFFFFFFFFFF; assign b = 64'h79DFFFFFFFFFFFFF;

    #10 $display("\n2**98 * 2**925:");
    #10 assign a = 64'h4610000000000000; assign b = 64'h79C0000000000000;
    #10 assign a = 64'h461FFFFFFFFFFFFF; assign b = 64'h79CFFFFFFFFFFFFF;

    #10 $display("\n2**99 * 2**924:");
    #10 assign a = 64'h4620000000000000; assign b = 64'h79B0000000000000;
    #10 assign a = 64'h462FFFFFFFFFFFFF; assign b = 64'h79BFFFFFFFFFFFFF;

    #10 $display("\n2**100 * 2**923:");
    #10 assign a = 64'h4630000000000000; assign b = 64'h79A0000000000000;
    #10 assign a = 64'h463FFFFFFFFFFFFF; assign b = 64'h79AFFFFFFFFFFFFF;

    #10 $display("\n2**101 * 2**922:");
    #10 assign a = 64'h4640000000000000; assign b = 64'h7990000000000000;
    #10 assign a = 64'h464FFFFFFFFFFFFF; assign b = 64'h799FFFFFFFFFFFFF;

    #10 $display("\n2**102 * 2**921:");
    #10 assign a = 64'h4650000000000000; assign b = 64'h7980000000000000;
    #10 assign a = 64'h465FFFFFFFFFFFFF; assign b = 64'h798FFFFFFFFFFFFF;

    #10 $display("\n2**103 * 2**920:");
    #10 assign a = 64'h4660000000000000; assign b = 64'h7970000000000000;
    #10 assign a = 64'h466FFFFFFFFFFFFF; assign b = 64'h797FFFFFFFFFFFFF;

    #10 $display("\n2**104 * 2**919:");
    #10 assign a = 64'h4670000000000000; assign b = 64'h7960000000000000;
    #10 assign a = 64'h467FFFFFFFFFFFFF; assign b = 64'h796FFFFFFFFFFFFF;

    #10 $display("\n2**105 * 2**918:");
    #10 assign a = 64'h4680000000000000; assign b = 64'h7950000000000000;
    #10 assign a = 64'h468FFFFFFFFFFFFF; assign b = 64'h795FFFFFFFFFFFFF;

    #10 $display("\n2**106 * 2**917:");
    #10 assign a = 64'h4690000000000000; assign b = 64'h7940000000000000;
    #10 assign a = 64'h469FFFFFFFFFFFFF; assign b = 64'h794FFFFFFFFFFFFF;

    #10 $display("\n2**107 * 2**916:");
    #10 assign a = 64'h46A0000000000000; assign b = 64'h7930000000000000;
    #10 assign a = 64'h46AFFFFFFFFFFFFF; assign b = 64'h793FFFFFFFFFFFFF;

    #10 $display("\n2**108 * 2**915:");
    #10 assign a = 64'h46B0000000000000; assign b = 64'h7920000000000000;
    #10 assign a = 64'h46BFFFFFFFFFFFFF; assign b = 64'h792FFFFFFFFFFFFF;

    #10 $display("\n2**109 * 2**914:");
    #10 assign a = 64'h46C0000000000000; assign b = 64'h7910000000000000;
    #10 assign a = 64'h46CFFFFFFFFFFFFF; assign b = 64'h791FFFFFFFFFFFFF;

    #10 $display("\n2**110 * 2**913:");
    #10 assign a = 64'h46D0000000000000; assign b = 64'h7900000000000000;
    #10 assign a = 64'h46DFFFFFFFFFFFFF; assign b = 64'h790FFFFFFFFFFFFF;

    #10 $display("\n2**111 * 2**912:");
    #10 assign a = 64'h46E0000000000000; assign b = 64'h78F0000000000000;
    #10 assign a = 64'h46EFFFFFFFFFFFFF; assign b = 64'h78FFFFFFFFFFFFFF;

    #10 $display("\n2**112 * 2**911:");
    #10 assign a = 64'h46F0000000000000; assign b = 64'h78E0000000000000;
    #10 assign a = 64'h46FFFFFFFFFFFFFF; assign b = 64'h78EFFFFFFFFFFFFF;

    #10 $display("\n2**113 * 2**910:");
    #10 assign a = 64'h4700000000000000; assign b = 64'h78D0000000000000;
    #10 assign a = 64'h470FFFFFFFFFFFFF; assign b = 64'h78DFFFFFFFFFFFFF;

    #10 $display("\n2**114 * 2**909:");
    #10 assign a = 64'h4710000000000000; assign b = 64'h78C0000000000000;
    #10 assign a = 64'h471FFFFFFFFFFFFF; assign b = 64'h78CFFFFFFFFFFFFF;

    #10 $display("\n2**115 * 2**908:");
    #10 assign a = 64'h4720000000000000; assign b = 64'h78B0000000000000;
    #10 assign a = 64'h472FFFFFFFFFFFFF; assign b = 64'h78BFFFFFFFFFFFFF;

    #10 $display("\n2**116 * 2**907:");
    #10 assign a = 64'h4730000000000000; assign b = 64'h78A0000000000000;
    #10 assign a = 64'h473FFFFFFFFFFFFF; assign b = 64'h78AFFFFFFFFFFFFF;

    #10 $display("\n2**117 * 2**906:");
    #10 assign a = 64'h4740000000000000; assign b = 64'h7890000000000000;
    #10 assign a = 64'h474FFFFFFFFFFFFF; assign b = 64'h789FFFFFFFFFFFFF;

    #10 $display("\n2**118 * 2**905:");
    #10 assign a = 64'h4750000000000000; assign b = 64'h7880000000000000;
    #10 assign a = 64'h475FFFFFFFFFFFFF; assign b = 64'h788FFFFFFFFFFFFF;

    #10 $display("\n2**119 * 2**904:");
    #10 assign a = 64'h4760000000000000; assign b = 64'h7870000000000000;
    #10 assign a = 64'h476FFFFFFFFFFFFF; assign b = 64'h787FFFFFFFFFFFFF;

    #10 $display("\n2**120 * 2**903:");
    #10 assign a = 64'h4770000000000000; assign b = 64'h7860000000000000;
    #10 assign a = 64'h477FFFFFFFFFFFFF; assign b = 64'h786FFFFFFFFFFFFF;

    #10 $display("\n2**121 * 2**902:");
    #10 assign a = 64'h4780000000000000; assign b = 64'h7850000000000000;
    #10 assign a = 64'h478FFFFFFFFFFFFF; assign b = 64'h785FFFFFFFFFFFFF;

    #10 $display("\n2**122 * 2**901:");
    #10 assign a = 64'h4790000000000000; assign b = 64'h7840000000000000;
    #10 assign a = 64'h479FFFFFFFFFFFFF; assign b = 64'h784FFFFFFFFFFFFF;

    #10 $display("\n2**123 * 2**900:");
    #10 assign a = 64'h47A0000000000000; assign b = 64'h7830000000000000;
    #10 assign a = 64'h47AFFFFFFFFFFFFF; assign b = 64'h783FFFFFFFFFFFFF;

    #10 $display("\n2**124 * 2**899:");
    #10 assign a = 64'h47B0000000000000; assign b = 64'h7820000000000000;
    #10 assign a = 64'h47BFFFFFFFFFFFFF; assign b = 64'h782FFFFFFFFFFFFF;

    #10 $display("\n2**125 * 2**898:");
    #10 assign a = 64'h47C0000000000000; assign b = 64'h7810000000000000;
    #10 assign a = 64'h47CFFFFFFFFFFFFF; assign b = 64'h781FFFFFFFFFFFFF;

    #10 $display("\n2**126 * 2**897:");
    #10 assign a = 64'h47D0000000000000; assign b = 64'h7800000000000000;
    #10 assign a = 64'h47DFFFFFFFFFFFFF; assign b = 64'h780FFFFFFFFFFFFF;

    #10 $display("\n2**127 * 2**896:");
    #10 assign a = 64'h47E0000000000000; assign b = 64'h77F0000000000000;
    #10 assign a = 64'h47EFFFFFFFFFFFFF; assign b = 64'h77FFFFFFFFFFFFFF;

    #10 $display("\n2**128 * 2**895:");
    #10 assign a = 64'h47F0000000000000; assign b = 64'h77E0000000000000;
    #10 assign a = 64'h47FFFFFFFFFFFFFF; assign b = 64'h77EFFFFFFFFFFFFF;

    #10 $display("\n2**129 * 2**894:");
    #10 assign a = 64'h4800000000000000; assign b = 64'h77D0000000000000;
    #10 assign a = 64'h480FFFFFFFFFFFFF; assign b = 64'h77DFFFFFFFFFFFFF;

    #10 $display("\n2**130 * 2**893:");
    #10 assign a = 64'h4810000000000000; assign b = 64'h77C0000000000000;
    #10 assign a = 64'h481FFFFFFFFFFFFF; assign b = 64'h77CFFFFFFFFFFFFF;

    #10 $display("\n2**131 * 2**892:");
    #10 assign a = 64'h4820000000000000; assign b = 64'h77B0000000000000;
    #10 assign a = 64'h482FFFFFFFFFFFFF; assign b = 64'h77BFFFFFFFFFFFFF;

    #10 $display("\n2**132 * 2**891:");
    #10 assign a = 64'h4830000000000000; assign b = 64'h77A0000000000000;
    #10 assign a = 64'h483FFFFFFFFFFFFF; assign b = 64'h77AFFFFFFFFFFFFF;

    #10 $display("\n2**133 * 2**890:");
    #10 assign a = 64'h4840000000000000; assign b = 64'h7790000000000000;
    #10 assign a = 64'h484FFFFFFFFFFFFF; assign b = 64'h779FFFFFFFFFFFFF;

    #10 $display("\n2**134 * 2**889:");
    #10 assign a = 64'h4850000000000000; assign b = 64'h7780000000000000;
    #10 assign a = 64'h485FFFFFFFFFFFFF; assign b = 64'h778FFFFFFFFFFFFF;

    #10 $display("\n2**135 * 2**888:");
    #10 assign a = 64'h4860000000000000; assign b = 64'h7770000000000000;
    #10 assign a = 64'h486FFFFFFFFFFFFF; assign b = 64'h777FFFFFFFFFFFFF;

    #10 $display("\n2**136 * 2**887:");
    #10 assign a = 64'h4870000000000000; assign b = 64'h7760000000000000;
    #10 assign a = 64'h487FFFFFFFFFFFFF; assign b = 64'h776FFFFFFFFFFFFF;

    #10 $display("\n2**137 * 2**886:");
    #10 assign a = 64'h4880000000000000; assign b = 64'h7750000000000000;
    #10 assign a = 64'h488FFFFFFFFFFFFF; assign b = 64'h775FFFFFFFFFFFFF;

    #10 $display("\n2**138 * 2**885:");
    #10 assign a = 64'h4890000000000000; assign b = 64'h7740000000000000;
    #10 assign a = 64'h489FFFFFFFFFFFFF; assign b = 64'h774FFFFFFFFFFFFF;

    #10 $display("\n2**139 * 2**884:");
    #10 assign a = 64'h48A0000000000000; assign b = 64'h7730000000000000;
    #10 assign a = 64'h48AFFFFFFFFFFFFF; assign b = 64'h773FFFFFFFFFFFFF;

    #10 $display("\n2**140 * 2**883:");
    #10 assign a = 64'h48B0000000000000; assign b = 64'h7720000000000000;
    #10 assign a = 64'h48BFFFFFFFFFFFFF; assign b = 64'h772FFFFFFFFFFFFF;

    #10 $display("\n2**141 * 2**882:");
    #10 assign a = 64'h48C0000000000000; assign b = 64'h7710000000000000;
    #10 assign a = 64'h48CFFFFFFFFFFFFF; assign b = 64'h771FFFFFFFFFFFFF;

    #10 $display("\n2**142 * 2**881:");
    #10 assign a = 64'h48D0000000000000; assign b = 64'h7700000000000000;
    #10 assign a = 64'h48DFFFFFFFFFFFFF; assign b = 64'h770FFFFFFFFFFFFF;

    #10 $display("\n2**143 * 2**880:");
    #10 assign a = 64'h48E0000000000000; assign b = 64'h76F0000000000000;
    #10 assign a = 64'h48EFFFFFFFFFFFFF; assign b = 64'h76FFFFFFFFFFFFFF;

    #10 $display("\n2**144 * 2**879:");
    #10 assign a = 64'h48F0000000000000; assign b = 64'h76E0000000000000;
    #10 assign a = 64'h48FFFFFFFFFFFFFF; assign b = 64'h76EFFFFFFFFFFFFF;

    #10 $display("\n2**145 * 2**878:");
    #10 assign a = 64'h4900000000000000; assign b = 64'h76D0000000000000;
    #10 assign a = 64'h490FFFFFFFFFFFFF; assign b = 64'h76DFFFFFFFFFFFFF;

    #10 $display("\n2**146 * 2**877:");
    #10 assign a = 64'h4910000000000000; assign b = 64'h76C0000000000000;
    #10 assign a = 64'h491FFFFFFFFFFFFF; assign b = 64'h76CFFFFFFFFFFFFF;

    #10 $display("\n2**147 * 2**876:");
    #10 assign a = 64'h4920000000000000; assign b = 64'h76B0000000000000;
    #10 assign a = 64'h492FFFFFFFFFFFFF; assign b = 64'h76BFFFFFFFFFFFFF;

    #10 $display("\n2**148 * 2**875:");
    #10 assign a = 64'h4930000000000000; assign b = 64'h76A0000000000000;
    #10 assign a = 64'h493FFFFFFFFFFFFF; assign b = 64'h76AFFFFFFFFFFFFF;

    #10 $display("\n2**149 * 2**874:");
    #10 assign a = 64'h4940000000000000; assign b = 64'h7690000000000000;
    #10 assign a = 64'h494FFFFFFFFFFFFF; assign b = 64'h769FFFFFFFFFFFFF;

    #10 $display("\n2**150 * 2**873:");
    #10 assign a = 64'h4950000000000000; assign b = 64'h7680000000000000;
    #10 assign a = 64'h495FFFFFFFFFFFFF; assign b = 64'h768FFFFFFFFFFFFF;

    #10 $display("\n2**151 * 2**872:");
    #10 assign a = 64'h4960000000000000; assign b = 64'h7670000000000000;
    #10 assign a = 64'h496FFFFFFFFFFFFF; assign b = 64'h767FFFFFFFFFFFFF;

    #10 $display("\n2**152 * 2**871:");
    #10 assign a = 64'h4970000000000000; assign b = 64'h7660000000000000;
    #10 assign a = 64'h497FFFFFFFFFFFFF; assign b = 64'h766FFFFFFFFFFFFF;

    #10 $display("\n2**153 * 2**870:");
    #10 assign a = 64'h4980000000000000; assign b = 64'h7650000000000000;
    #10 assign a = 64'h498FFFFFFFFFFFFF; assign b = 64'h765FFFFFFFFFFFFF;

    #10 $display("\n2**154 * 2**869:");
    #10 assign a = 64'h4990000000000000; assign b = 64'h7640000000000000;
    #10 assign a = 64'h499FFFFFFFFFFFFF; assign b = 64'h764FFFFFFFFFFFFF;

    #10 $display("\n2**155 * 2**868:");
    #10 assign a = 64'h49A0000000000000; assign b = 64'h7630000000000000;
    #10 assign a = 64'h49AFFFFFFFFFFFFF; assign b = 64'h763FFFFFFFFFFFFF;

    #10 $display("\n2**156 * 2**867:");
    #10 assign a = 64'h49B0000000000000; assign b = 64'h7620000000000000;
    #10 assign a = 64'h49BFFFFFFFFFFFFF; assign b = 64'h762FFFFFFFFFFFFF;

    #10 $display("\n2**157 * 2**866:");
    #10 assign a = 64'h49C0000000000000; assign b = 64'h7610000000000000;
    #10 assign a = 64'h49CFFFFFFFFFFFFF; assign b = 64'h761FFFFFFFFFFFFF;

    #10 $display("\n2**158 * 2**865:");
    #10 assign a = 64'h49D0000000000000; assign b = 64'h7600000000000000;
    #10 assign a = 64'h49DFFFFFFFFFFFFF; assign b = 64'h760FFFFFFFFFFFFF;

    #10 $display("\n2**159 * 2**864:");
    #10 assign a = 64'h49E0000000000000; assign b = 64'h75F0000000000000;
    #10 assign a = 64'h49EFFFFFFFFFFFFF; assign b = 64'h75FFFFFFFFFFFFFF;

    #10 $display("\n2**160 * 2**863:");
    #10 assign a = 64'h49F0000000000000; assign b = 64'h75E0000000000000;
    #10 assign a = 64'h49FFFFFFFFFFFFFF; assign b = 64'h75EFFFFFFFFFFFFF;

    #10 $display("\n2**161 * 2**862:");
    #10 assign a = 64'h4A00000000000000; assign b = 64'h75D0000000000000;
    #10 assign a = 64'h4A0FFFFFFFFFFFFF; assign b = 64'h75DFFFFFFFFFFFFF;

    #10 $display("\n2**162 * 2**861:");
    #10 assign a = 64'h4A10000000000000; assign b = 64'h75C0000000000000;
    #10 assign a = 64'h4A1FFFFFFFFFFFFF; assign b = 64'h75CFFFFFFFFFFFFF;

    #10 $display("\n2**163 * 2**860:");
    #10 assign a = 64'h4A20000000000000; assign b = 64'h75B0000000000000;
    #10 assign a = 64'h4A2FFFFFFFFFFFFF; assign b = 64'h75BFFFFFFFFFFFFF;

    #10 $display("\n2**164 * 2**859:");
    #10 assign a = 64'h4A30000000000000; assign b = 64'h75A0000000000000;
    #10 assign a = 64'h4A3FFFFFFFFFFFFF; assign b = 64'h75AFFFFFFFFFFFFF;

    #10 $display("\n2**165 * 2**858:");
    #10 assign a = 64'h4A40000000000000; assign b = 64'h7590000000000000;
    #10 assign a = 64'h4A4FFFFFFFFFFFFF; assign b = 64'h759FFFFFFFFFFFFF;

    #10 $display("\n2**166 * 2**857:");
    #10 assign a = 64'h4A50000000000000; assign b = 64'h7580000000000000;
    #10 assign a = 64'h4A5FFFFFFFFFFFFF; assign b = 64'h758FFFFFFFFFFFFF;

    #10 $display("\n2**167 * 2**856:");
    #10 assign a = 64'h4A60000000000000; assign b = 64'h7570000000000000;
    #10 assign a = 64'h4A6FFFFFFFFFFFFF; assign b = 64'h757FFFFFFFFFFFFF;

    #10 $display("\n2**168 * 2**855:");
    #10 assign a = 64'h4A70000000000000; assign b = 64'h7560000000000000;
    #10 assign a = 64'h4A7FFFFFFFFFFFFF; assign b = 64'h756FFFFFFFFFFFFF;

    #10 $display("\n2**169 * 2**854:");
    #10 assign a = 64'h4A80000000000000; assign b = 64'h7550000000000000;
    #10 assign a = 64'h4A8FFFFFFFFFFFFF; assign b = 64'h755FFFFFFFFFFFFF;

    #10 $display("\n2**170 * 2**853:");
    #10 assign a = 64'h4A90000000000000; assign b = 64'h7540000000000000;
    #10 assign a = 64'h4A9FFFFFFFFFFFFF; assign b = 64'h754FFFFFFFFFFFFF;

    #10 $display("\n2**171 * 2**852:");
    #10 assign a = 64'h4AA0000000000000; assign b = 64'h7530000000000000;
    #10 assign a = 64'h4AAFFFFFFFFFFFFF; assign b = 64'h753FFFFFFFFFFFFF;

    #10 $display("\n2**172 * 2**851:");
    #10 assign a = 64'h4AB0000000000000; assign b = 64'h7520000000000000;
    #10 assign a = 64'h4ABFFFFFFFFFFFFF; assign b = 64'h752FFFFFFFFFFFFF;

    #10 $display("\n2**173 * 2**850:");
    #10 assign a = 64'h4AC0000000000000; assign b = 64'h7510000000000000;
    #10 assign a = 64'h4ACFFFFFFFFFFFFF; assign b = 64'h751FFFFFFFFFFFFF;

    #10 $display("\n2**174 * 2**849:");
    #10 assign a = 64'h4AD0000000000000; assign b = 64'h7500000000000000;
    #10 assign a = 64'h4ADFFFFFFFFFFFFF; assign b = 64'h750FFFFFFFFFFFFF;

    #10 $display("\n2**175 * 2**848:");
    #10 assign a = 64'h4AE0000000000000; assign b = 64'h74F0000000000000;
    #10 assign a = 64'h4AEFFFFFFFFFFFFF; assign b = 64'h74FFFFFFFFFFFFFF;

    #10 $display("\n2**176 * 2**847:");
    #10 assign a = 64'h4AF0000000000000; assign b = 64'h74E0000000000000;
    #10 assign a = 64'h4AFFFFFFFFFFFFFF; assign b = 64'h74EFFFFFFFFFFFFF;

    #10 $display("\n2**177 * 2**846:");
    #10 assign a = 64'h4B00000000000000; assign b = 64'h74D0000000000000;
    #10 assign a = 64'h4B0FFFFFFFFFFFFF; assign b = 64'h74DFFFFFFFFFFFFF;

    #10 $display("\n2**178 * 2**845:");
    #10 assign a = 64'h4B10000000000000; assign b = 64'h74C0000000000000;
    #10 assign a = 64'h4B1FFFFFFFFFFFFF; assign b = 64'h74CFFFFFFFFFFFFF;

    #10 $display("\n2**179 * 2**844:");
    #10 assign a = 64'h4B20000000000000; assign b = 64'h74B0000000000000;
    #10 assign a = 64'h4B2FFFFFFFFFFFFF; assign b = 64'h74BFFFFFFFFFFFFF;

    #10 $display("\n2**180 * 2**843:");
    #10 assign a = 64'h4B30000000000000; assign b = 64'h74A0000000000000;
    #10 assign a = 64'h4B3FFFFFFFFFFFFF; assign b = 64'h74AFFFFFFFFFFFFF;

    #10 $display("\n2**181 * 2**842:");
    #10 assign a = 64'h4B40000000000000; assign b = 64'h7490000000000000;
    #10 assign a = 64'h4B4FFFFFFFFFFFFF; assign b = 64'h749FFFFFFFFFFFFF;

    #10 $display("\n2**182 * 2**841:");
    #10 assign a = 64'h4B50000000000000; assign b = 64'h7480000000000000;
    #10 assign a = 64'h4B5FFFFFFFFFFFFF; assign b = 64'h748FFFFFFFFFFFFF;

    #10 $display("\n2**183 * 2**840:");
    #10 assign a = 64'h4B60000000000000; assign b = 64'h7470000000000000;
    #10 assign a = 64'h4B6FFFFFFFFFFFFF; assign b = 64'h747FFFFFFFFFFFFF;

    #10 $display("\n2**184 * 2**839:");
    #10 assign a = 64'h4B70000000000000; assign b = 64'h7460000000000000;
    #10 assign a = 64'h4B7FFFFFFFFFFFFF; assign b = 64'h746FFFFFFFFFFFFF;

    #10 $display("\n2**185 * 2**838:");
    #10 assign a = 64'h4B80000000000000; assign b = 64'h7450000000000000;
    #10 assign a = 64'h4B8FFFFFFFFFFFFF; assign b = 64'h745FFFFFFFFFFFFF;

    #10 $display("\n2**186 * 2**837:");
    #10 assign a = 64'h4B90000000000000; assign b = 64'h7440000000000000;
    #10 assign a = 64'h4B9FFFFFFFFFFFFF; assign b = 64'h744FFFFFFFFFFFFF;

    #10 $display("\n2**187 * 2**836:");
    #10 assign a = 64'h4BA0000000000000; assign b = 64'h7430000000000000;
    #10 assign a = 64'h4BAFFFFFFFFFFFFF; assign b = 64'h743FFFFFFFFFFFFF;

    #10 $display("\n2**188 * 2**835:");
    #10 assign a = 64'h4BB0000000000000; assign b = 64'h7420000000000000;
    #10 assign a = 64'h4BBFFFFFFFFFFFFF; assign b = 64'h742FFFFFFFFFFFFF;

    #10 $display("\n2**189 * 2**834:");
    #10 assign a = 64'h4BC0000000000000; assign b = 64'h7410000000000000;
    #10 assign a = 64'h4BCFFFFFFFFFFFFF; assign b = 64'h741FFFFFFFFFFFFF;

    #10 $display("\n2**190 * 2**833:");
    #10 assign a = 64'h4BD0000000000000; assign b = 64'h7400000000000000;
    #10 assign a = 64'h4BDFFFFFFFFFFFFF; assign b = 64'h740FFFFFFFFFFFFF;

    #10 $display("\n2**191 * 2**832:");
    #10 assign a = 64'h4BE0000000000000; assign b = 64'h73F0000000000000;
    #10 assign a = 64'h4BEFFFFFFFFFFFFF; assign b = 64'h73FFFFFFFFFFFFFF;

    #10 $display("\n2**192 * 2**831:");
    #10 assign a = 64'h4BF0000000000000; assign b = 64'h73E0000000000000;
    #10 assign a = 64'h4BFFFFFFFFFFFFFF; assign b = 64'h73EFFFFFFFFFFFFF;

    #10 $display("\n2**193 * 2**830:");
    #10 assign a = 64'h4C00000000000000; assign b = 64'h73D0000000000000;
    #10 assign a = 64'h4C0FFFFFFFFFFFFF; assign b = 64'h73DFFFFFFFFFFFFF;

    #10 $display("\n2**194 * 2**829:");
    #10 assign a = 64'h4C10000000000000; assign b = 64'h73C0000000000000;
    #10 assign a = 64'h4C1FFFFFFFFFFFFF; assign b = 64'h73CFFFFFFFFFFFFF;

    #10 $display("\n2**195 * 2**828:");
    #10 assign a = 64'h4C20000000000000; assign b = 64'h73B0000000000000;
    #10 assign a = 64'h4C2FFFFFFFFFFFFF; assign b = 64'h73BFFFFFFFFFFFFF;

    #10 $display("\n2**196 * 2**827:");
    #10 assign a = 64'h4C30000000000000; assign b = 64'h73A0000000000000;
    #10 assign a = 64'h4C3FFFFFFFFFFFFF; assign b = 64'h73AFFFFFFFFFFFFF;

    #10 $display("\n2**197 * 2**826:");
    #10 assign a = 64'h4C40000000000000; assign b = 64'h7390000000000000;
    #10 assign a = 64'h4C4FFFFFFFFFFFFF; assign b = 64'h739FFFFFFFFFFFFF;

    #10 $display("\n2**198 * 2**825:");
    #10 assign a = 64'h4C50000000000000; assign b = 64'h7380000000000000;
    #10 assign a = 64'h4C5FFFFFFFFFFFFF; assign b = 64'h738FFFFFFFFFFFFF;

    #10 $display("\n2**199 * 2**824:");
    #10 assign a = 64'h4C60000000000000; assign b = 64'h7370000000000000;
    #10 assign a = 64'h4C6FFFFFFFFFFFFF; assign b = 64'h737FFFFFFFFFFFFF;

    #10 $display("\n2**200 * 2**823:");
    #10 assign a = 64'h4C70000000000000; assign b = 64'h7360000000000000;
    #10 assign a = 64'h4C7FFFFFFFFFFFFF; assign b = 64'h736FFFFFFFFFFFFF;

    #10 $display("\n2**201 * 2**822:");
    #10 assign a = 64'h4C80000000000000; assign b = 64'h7350000000000000;
    #10 assign a = 64'h4C8FFFFFFFFFFFFF; assign b = 64'h735FFFFFFFFFFFFF;

    #10 $display("\n2**202 * 2**821:");
    #10 assign a = 64'h4C90000000000000; assign b = 64'h7340000000000000;
    #10 assign a = 64'h4C9FFFFFFFFFFFFF; assign b = 64'h734FFFFFFFFFFFFF;

    #10 $display("\n2**203 * 2**820:");
    #10 assign a = 64'h4CA0000000000000; assign b = 64'h7330000000000000;
    #10 assign a = 64'h4CAFFFFFFFFFFFFF; assign b = 64'h733FFFFFFFFFFFFF;

    #10 $display("\n2**204 * 2**819:");
    #10 assign a = 64'h4CB0000000000000; assign b = 64'h7320000000000000;
    #10 assign a = 64'h4CBFFFFFFFFFFFFF; assign b = 64'h732FFFFFFFFFFFFF;

    #10 $display("\n2**205 * 2**818:");
    #10 assign a = 64'h4CC0000000000000; assign b = 64'h7310000000000000;
    #10 assign a = 64'h4CCFFFFFFFFFFFFF; assign b = 64'h731FFFFFFFFFFFFF;

    #10 $display("\n2**206 * 2**817:");
    #10 assign a = 64'h4CD0000000000000; assign b = 64'h7300000000000000;
    #10 assign a = 64'h4CDFFFFFFFFFFFFF; assign b = 64'h730FFFFFFFFFFFFF;

    #10 $display("\n2**207 * 2**816:");
    #10 assign a = 64'h4CE0000000000000; assign b = 64'h72F0000000000000;
    #10 assign a = 64'h4CEFFFFFFFFFFFFF; assign b = 64'h72FFFFFFFFFFFFFF;

    #10 $display("\n2**208 * 2**815:");
    #10 assign a = 64'h4CF0000000000000; assign b = 64'h72E0000000000000;
    #10 assign a = 64'h4CFFFFFFFFFFFFFF; assign b = 64'h72EFFFFFFFFFFFFF;

    #10 $display("\n2**209 * 2**814:");
    #10 assign a = 64'h4D00000000000000; assign b = 64'h72D0000000000000;
    #10 assign a = 64'h4D0FFFFFFFFFFFFF; assign b = 64'h72DFFFFFFFFFFFFF;

    #10 $display("\n2**210 * 2**813:");
    #10 assign a = 64'h4D10000000000000; assign b = 64'h72C0000000000000;
    #10 assign a = 64'h4D1FFFFFFFFFFFFF; assign b = 64'h72CFFFFFFFFFFFFF;

    #10 $display("\n2**211 * 2**812:");
    #10 assign a = 64'h4D20000000000000; assign b = 64'h72B0000000000000;
    #10 assign a = 64'h4D2FFFFFFFFFFFFF; assign b = 64'h72BFFFFFFFFFFFFF;

    #10 $display("\n2**212 * 2**811:");
    #10 assign a = 64'h4D30000000000000; assign b = 64'h72A0000000000000;
    #10 assign a = 64'h4D3FFFFFFFFFFFFF; assign b = 64'h72AFFFFFFFFFFFFF;

    #10 $display("\n2**213 * 2**810:");
    #10 assign a = 64'h4D40000000000000; assign b = 64'h7290000000000000;
    #10 assign a = 64'h4D4FFFFFFFFFFFFF; assign b = 64'h729FFFFFFFFFFFFF;

    #10 $display("\n2**214 * 2**809:");
    #10 assign a = 64'h4D50000000000000; assign b = 64'h7280000000000000;
    #10 assign a = 64'h4D5FFFFFFFFFFFFF; assign b = 64'h728FFFFFFFFFFFFF;

    #10 $display("\n2**215 * 2**808:");
    #10 assign a = 64'h4D60000000000000; assign b = 64'h7270000000000000;
    #10 assign a = 64'h4D6FFFFFFFFFFFFF; assign b = 64'h727FFFFFFFFFFFFF;

    #10 $display("\n2**216 * 2**807:");
    #10 assign a = 64'h4D70000000000000; assign b = 64'h7260000000000000;
    #10 assign a = 64'h4D7FFFFFFFFFFFFF; assign b = 64'h726FFFFFFFFFFFFF;

    #10 $display("\n2**217 * 2**806:");
    #10 assign a = 64'h4D80000000000000; assign b = 64'h7250000000000000;
    #10 assign a = 64'h4D8FFFFFFFFFFFFF; assign b = 64'h725FFFFFFFFFFFFF;

    #10 $display("\n2**218 * 2**805:");
    #10 assign a = 64'h4D90000000000000; assign b = 64'h7240000000000000;
    #10 assign a = 64'h4D9FFFFFFFFFFFFF; assign b = 64'h724FFFFFFFFFFFFF;

    #10 $display("\n2**219 * 2**804:");
    #10 assign a = 64'h4DA0000000000000; assign b = 64'h7230000000000000;
    #10 assign a = 64'h4DAFFFFFFFFFFFFF; assign b = 64'h723FFFFFFFFFFFFF;

    #10 $display("\n2**220 * 2**803:");
    #10 assign a = 64'h4DB0000000000000; assign b = 64'h7220000000000000;
    #10 assign a = 64'h4DBFFFFFFFFFFFFF; assign b = 64'h722FFFFFFFFFFFFF;

    #10 $display("\n2**221 * 2**802:");
    #10 assign a = 64'h4DC0000000000000; assign b = 64'h7210000000000000;
    #10 assign a = 64'h4DCFFFFFFFFFFFFF; assign b = 64'h721FFFFFFFFFFFFF;

    #10 $display("\n2**222 * 2**801:");
    #10 assign a = 64'h4DD0000000000000; assign b = 64'h7200000000000000;
    #10 assign a = 64'h4DDFFFFFFFFFFFFF; assign b = 64'h720FFFFFFFFFFFFF;

    #10 $display("\n2**223 * 2**800:");
    #10 assign a = 64'h4DE0000000000000; assign b = 64'h71F0000000000000;
    #10 assign a = 64'h4DEFFFFFFFFFFFFF; assign b = 64'h71FFFFFFFFFFFFFF;

    #10 $display("\n2**224 * 2**799:");
    #10 assign a = 64'h4DF0000000000000; assign b = 64'h71E0000000000000;
    #10 assign a = 64'h4DFFFFFFFFFFFFFF; assign b = 64'h71EFFFFFFFFFFFFF;

    #10 $display("\n2**225 * 2**798:");
    #10 assign a = 64'h4E00000000000000; assign b = 64'h71D0000000000000;
    #10 assign a = 64'h4E0FFFFFFFFFFFFF; assign b = 64'h71DFFFFFFFFFFFFF;

    #10 $display("\n2**226 * 2**797:");
    #10 assign a = 64'h4E10000000000000; assign b = 64'h71C0000000000000;
    #10 assign a = 64'h4E1FFFFFFFFFFFFF; assign b = 64'h71CFFFFFFFFFFFFF;

    #10 $display("\n2**227 * 2**796:");
    #10 assign a = 64'h4E20000000000000; assign b = 64'h71B0000000000000;
    #10 assign a = 64'h4E2FFFFFFFFFFFFF; assign b = 64'h71BFFFFFFFFFFFFF;

    #10 $display("\n2**228 * 2**795:");
    #10 assign a = 64'h4E30000000000000; assign b = 64'h71A0000000000000;
    #10 assign a = 64'h4E3FFFFFFFFFFFFF; assign b = 64'h71AFFFFFFFFFFFFF;

    #10 $display("\n2**229 * 2**794:");
    #10 assign a = 64'h4E40000000000000; assign b = 64'h7190000000000000;
    #10 assign a = 64'h4E4FFFFFFFFFFFFF; assign b = 64'h719FFFFFFFFFFFFF;

    #10 $display("\n2**230 * 2**793:");
    #10 assign a = 64'h4E50000000000000; assign b = 64'h7180000000000000;
    #10 assign a = 64'h4E5FFFFFFFFFFFFF; assign b = 64'h718FFFFFFFFFFFFF;

    #10 $display("\n2**231 * 2**792:");
    #10 assign a = 64'h4E60000000000000; assign b = 64'h7170000000000000;
    #10 assign a = 64'h4E6FFFFFFFFFFFFF; assign b = 64'h717FFFFFFFFFFFFF;

    #10 $display("\n2**232 * 2**791:");
    #10 assign a = 64'h4E70000000000000; assign b = 64'h7160000000000000;
    #10 assign a = 64'h4E7FFFFFFFFFFFFF; assign b = 64'h716FFFFFFFFFFFFF;

    #10 $display("\n2**233 * 2**790:");
    #10 assign a = 64'h4E80000000000000; assign b = 64'h7150000000000000;
    #10 assign a = 64'h4E8FFFFFFFFFFFFF; assign b = 64'h715FFFFFFFFFFFFF;

    #10 $display("\n2**234 * 2**789:");
    #10 assign a = 64'h4E90000000000000; assign b = 64'h7140000000000000;
    #10 assign a = 64'h4E9FFFFFFFFFFFFF; assign b = 64'h714FFFFFFFFFFFFF;

    #10 $display("\n2**235 * 2**788:");
    #10 assign a = 64'h4EA0000000000000; assign b = 64'h7130000000000000;
    #10 assign a = 64'h4EAFFFFFFFFFFFFF; assign b = 64'h713FFFFFFFFFFFFF;

    #10 $display("\n2**236 * 2**787:");
    #10 assign a = 64'h4EB0000000000000; assign b = 64'h7120000000000000;
    #10 assign a = 64'h4EBFFFFFFFFFFFFF; assign b = 64'h712FFFFFFFFFFFFF;

    #10 $display("\n2**237 * 2**786:");
    #10 assign a = 64'h4EC0000000000000; assign b = 64'h7110000000000000;
    #10 assign a = 64'h4ECFFFFFFFFFFFFF; assign b = 64'h711FFFFFFFFFFFFF;

    #10 $display("\n2**238 * 2**785:");
    #10 assign a = 64'h4ED0000000000000; assign b = 64'h7100000000000000;
    #10 assign a = 64'h4EDFFFFFFFFFFFFF; assign b = 64'h710FFFFFFFFFFFFF;

    #10 $display("\n2**239 * 2**784:");
    #10 assign a = 64'h4EE0000000000000; assign b = 64'h70F0000000000000;
    #10 assign a = 64'h4EEFFFFFFFFFFFFF; assign b = 64'h70FFFFFFFFFFFFFF;

    #10 $display("\n2**240 * 2**783:");
    #10 assign a = 64'h4EF0000000000000; assign b = 64'h70E0000000000000;
    #10 assign a = 64'h4EFFFFFFFFFFFFFF; assign b = 64'h70EFFFFFFFFFFFFF;

    #10 $display("\n2**241 * 2**782:");
    #10 assign a = 64'h4F00000000000000; assign b = 64'h70D0000000000000;
    #10 assign a = 64'h4F0FFFFFFFFFFFFF; assign b = 64'h70DFFFFFFFFFFFFF;

    #10 $display("\n2**242 * 2**781:");
    #10 assign a = 64'h4F10000000000000; assign b = 64'h70C0000000000000;
    #10 assign a = 64'h4F1FFFFFFFFFFFFF; assign b = 64'h70CFFFFFFFFFFFFF;

    #10 $display("\n2**243 * 2**780:");
    #10 assign a = 64'h4F20000000000000; assign b = 64'h70B0000000000000;
    #10 assign a = 64'h4F2FFFFFFFFFFFFF; assign b = 64'h70BFFFFFFFFFFFFF;

    #10 $display("\n2**244 * 2**779:");
    #10 assign a = 64'h4F30000000000000; assign b = 64'h70A0000000000000;
    #10 assign a = 64'h4F3FFFFFFFFFFFFF; assign b = 64'h70AFFFFFFFFFFFFF;

    #10 $display("\n2**245 * 2**778:");
    #10 assign a = 64'h4F40000000000000; assign b = 64'h7090000000000000;
    #10 assign a = 64'h4F4FFFFFFFFFFFFF; assign b = 64'h709FFFFFFFFFFFFF;

    #10 $display("\n2**246 * 2**777:");
    #10 assign a = 64'h4F50000000000000; assign b = 64'h7080000000000000;
    #10 assign a = 64'h4F5FFFFFFFFFFFFF; assign b = 64'h708FFFFFFFFFFFFF;

    #10 $display("\n2**247 * 2**776:");
    #10 assign a = 64'h4F60000000000000; assign b = 64'h7070000000000000;
    #10 assign a = 64'h4F6FFFFFFFFFFFFF; assign b = 64'h707FFFFFFFFFFFFF;

    #10 $display("\n2**248 * 2**775:");
    #10 assign a = 64'h4F70000000000000; assign b = 64'h7060000000000000;
    #10 assign a = 64'h4F7FFFFFFFFFFFFF; assign b = 64'h706FFFFFFFFFFFFF;

    #10 $display("\n2**249 * 2**774:");
    #10 assign a = 64'h4F80000000000000; assign b = 64'h7050000000000000;
    #10 assign a = 64'h4F8FFFFFFFFFFFFF; assign b = 64'h705FFFFFFFFFFFFF;

    #10 $display("\n2**250 * 2**773:");
    #10 assign a = 64'h4F90000000000000; assign b = 64'h7040000000000000;
    #10 assign a = 64'h4F9FFFFFFFFFFFFF; assign b = 64'h704FFFFFFFFFFFFF;

    #10 $display("\n2**251 * 2**772:");
    #10 assign a = 64'h4FA0000000000000; assign b = 64'h7030000000000000;
    #10 assign a = 64'h4FAFFFFFFFFFFFFF; assign b = 64'h703FFFFFFFFFFFFF;

    #10 $display("\n2**252 * 2**771:");
    #10 assign a = 64'h4FB0000000000000; assign b = 64'h7020000000000000;
    #10 assign a = 64'h4FBFFFFFFFFFFFFF; assign b = 64'h702FFFFFFFFFFFFF;

    #10 $display("\n2**253 * 2**770:");
    #10 assign a = 64'h4FC0000000000000; assign b = 64'h7010000000000000;
    #10 assign a = 64'h4FCFFFFFFFFFFFFF; assign b = 64'h701FFFFFFFFFFFFF;

    #10 $display("\n2**254 * 2**769:");
    #10 assign a = 64'h4FD0000000000000; assign b = 64'h7000000000000000;
    #10 assign a = 64'h4FDFFFFFFFFFFFFF; assign b = 64'h700FFFFFFFFFFFFF;

    #10 $display("\n2**255 * 2**768:");
    #10 assign a = 64'h4FE0000000000000; assign b = 64'h6FF0000000000000;
    #10 assign a = 64'h4FEFFFFFFFFFFFFF; assign b = 64'h6FFFFFFFFFFFFFFF;

    #10 $display("\n2**256 * 2**767:");
    #10 assign a = 64'h4FF0000000000000; assign b = 64'h6FE0000000000000;
    #10 assign a = 64'h4FFFFFFFFFFFFFFF; assign b = 64'h6FEFFFFFFFFFFFFF;

    #10 $display("\n2**257 * 2**766:");
    #10 assign a = 64'h5000000000000000; assign b = 64'h6FD0000000000000;
    #10 assign a = 64'h500FFFFFFFFFFFFF; assign b = 64'h6FDFFFFFFFFFFFFF;

    #10 $display("\n2**258 * 2**765:");
    #10 assign a = 64'h5010000000000000; assign b = 64'h6FC0000000000000;
    #10 assign a = 64'h501FFFFFFFFFFFFF; assign b = 64'h6FCFFFFFFFFFFFFF;

    #10 $display("\n2**259 * 2**764:");
    #10 assign a = 64'h5020000000000000; assign b = 64'h6FB0000000000000;
    #10 assign a = 64'h502FFFFFFFFFFFFF; assign b = 64'h6FBFFFFFFFFFFFFF;

    #10 $display("\n2**260 * 2**763:");
    #10 assign a = 64'h5030000000000000; assign b = 64'h6FA0000000000000;
    #10 assign a = 64'h503FFFFFFFFFFFFF; assign b = 64'h6FAFFFFFFFFFFFFF;

    #10 $display("\n2**261 * 2**762:");
    #10 assign a = 64'h5040000000000000; assign b = 64'h6F90000000000000;
    #10 assign a = 64'h504FFFFFFFFFFFFF; assign b = 64'h6F9FFFFFFFFFFFFF;

    #10 $display("\n2**262 * 2**761:");
    #10 assign a = 64'h5050000000000000; assign b = 64'h6F80000000000000;
    #10 assign a = 64'h505FFFFFFFFFFFFF; assign b = 64'h6F8FFFFFFFFFFFFF;

    #10 $display("\n2**263 * 2**760:");
    #10 assign a = 64'h5060000000000000; assign b = 64'h6F70000000000000;
    #10 assign a = 64'h506FFFFFFFFFFFFF; assign b = 64'h6F7FFFFFFFFFFFFF;

    #10 $display("\n2**264 * 2**759:");
    #10 assign a = 64'h5070000000000000; assign b = 64'h6F60000000000000;
    #10 assign a = 64'h507FFFFFFFFFFFFF; assign b = 64'h6F6FFFFFFFFFFFFF;

    #10 $display("\n2**265 * 2**758:");
    #10 assign a = 64'h5080000000000000; assign b = 64'h6F50000000000000;
    #10 assign a = 64'h508FFFFFFFFFFFFF; assign b = 64'h6F5FFFFFFFFFFFFF;

    #10 $display("\n2**266 * 2**757:");
    #10 assign a = 64'h5090000000000000; assign b = 64'h6F40000000000000;
    #10 assign a = 64'h509FFFFFFFFFFFFF; assign b = 64'h6F4FFFFFFFFFFFFF;

    #10 $display("\n2**267 * 2**756:");
    #10 assign a = 64'h50A0000000000000; assign b = 64'h6F30000000000000;
    #10 assign a = 64'h50AFFFFFFFFFFFFF; assign b = 64'h6F3FFFFFFFFFFFFF;

    #10 $display("\n2**268 * 2**755:");
    #10 assign a = 64'h50B0000000000000; assign b = 64'h6F20000000000000;
    #10 assign a = 64'h50BFFFFFFFFFFFFF; assign b = 64'h6F2FFFFFFFFFFFFF;

    #10 $display("\n2**269 * 2**754:");
    #10 assign a = 64'h50C0000000000000; assign b = 64'h6F10000000000000;
    #10 assign a = 64'h50CFFFFFFFFFFFFF; assign b = 64'h6F1FFFFFFFFFFFFF;

    #10 $display("\n2**270 * 2**753:");
    #10 assign a = 64'h50D0000000000000; assign b = 64'h6F00000000000000;
    #10 assign a = 64'h50DFFFFFFFFFFFFF; assign b = 64'h6F0FFFFFFFFFFFFF;

    #10 $display("\n2**271 * 2**752:");
    #10 assign a = 64'h50E0000000000000; assign b = 64'h6EF0000000000000;
    #10 assign a = 64'h50EFFFFFFFFFFFFF; assign b = 64'h6EFFFFFFFFFFFFFF;

    #10 $display("\n2**272 * 2**751:");
    #10 assign a = 64'h50F0000000000000; assign b = 64'h6EE0000000000000;
    #10 assign a = 64'h50FFFFFFFFFFFFFF; assign b = 64'h6EEFFFFFFFFFFFFF;

    #10 $display("\n2**273 * 2**750:");
    #10 assign a = 64'h5100000000000000; assign b = 64'h6ED0000000000000;
    #10 assign a = 64'h510FFFFFFFFFFFFF; assign b = 64'h6EDFFFFFFFFFFFFF;

    #10 $display("\n2**274 * 2**749:");
    #10 assign a = 64'h5110000000000000; assign b = 64'h6EC0000000000000;
    #10 assign a = 64'h511FFFFFFFFFFFFF; assign b = 64'h6ECFFFFFFFFFFFFF;

    #10 $display("\n2**275 * 2**748:");
    #10 assign a = 64'h5120000000000000; assign b = 64'h6EB0000000000000;
    #10 assign a = 64'h512FFFFFFFFFFFFF; assign b = 64'h6EBFFFFFFFFFFFFF;

    #10 $display("\n2**276 * 2**747:");
    #10 assign a = 64'h5130000000000000; assign b = 64'h6EA0000000000000;
    #10 assign a = 64'h513FFFFFFFFFFFFF; assign b = 64'h6EAFFFFFFFFFFFFF;

    #10 $display("\n2**277 * 2**746:");
    #10 assign a = 64'h5140000000000000; assign b = 64'h6E90000000000000;
    #10 assign a = 64'h514FFFFFFFFFFFFF; assign b = 64'h6E9FFFFFFFFFFFFF;

    #10 $display("\n2**278 * 2**745:");
    #10 assign a = 64'h5150000000000000; assign b = 64'h6E80000000000000;
    #10 assign a = 64'h515FFFFFFFFFFFFF; assign b = 64'h6E8FFFFFFFFFFFFF;

    #10 $display("\n2**279 * 2**744:");
    #10 assign a = 64'h5160000000000000; assign b = 64'h6E70000000000000;
    #10 assign a = 64'h516FFFFFFFFFFFFF; assign b = 64'h6E7FFFFFFFFFFFFF;

    #10 $display("\n2**280 * 2**743:");
    #10 assign a = 64'h5170000000000000; assign b = 64'h6E60000000000000;
    #10 assign a = 64'h517FFFFFFFFFFFFF; assign b = 64'h6E6FFFFFFFFFFFFF;

    #10 $display("\n2**281 * 2**742:");
    #10 assign a = 64'h5180000000000000; assign b = 64'h6E50000000000000;
    #10 assign a = 64'h518FFFFFFFFFFFFF; assign b = 64'h6E5FFFFFFFFFFFFF;

    #10 $display("\n2**282 * 2**741:");
    #10 assign a = 64'h5190000000000000; assign b = 64'h6E40000000000000;
    #10 assign a = 64'h519FFFFFFFFFFFFF; assign b = 64'h6E4FFFFFFFFFFFFF;

    #10 $display("\n2**283 * 2**740:");
    #10 assign a = 64'h51A0000000000000; assign b = 64'h6E30000000000000;
    #10 assign a = 64'h51AFFFFFFFFFFFFF; assign b = 64'h6E3FFFFFFFFFFFFF;

    #10 $display("\n2**284 * 2**739:");
    #10 assign a = 64'h51B0000000000000; assign b = 64'h6E20000000000000;
    #10 assign a = 64'h51BFFFFFFFFFFFFF; assign b = 64'h6E2FFFFFFFFFFFFF;

    #10 $display("\n2**285 * 2**738:");
    #10 assign a = 64'h51C0000000000000; assign b = 64'h6E10000000000000;
    #10 assign a = 64'h51CFFFFFFFFFFFFF; assign b = 64'h6E1FFFFFFFFFFFFF;

    #10 $display("\n2**286 * 2**737:");
    #10 assign a = 64'h51D0000000000000; assign b = 64'h6E00000000000000;
    #10 assign a = 64'h51DFFFFFFFFFFFFF; assign b = 64'h6E0FFFFFFFFFFFFF;

    #10 $display("\n2**287 * 2**736:");
    #10 assign a = 64'h51E0000000000000; assign b = 64'h6DF0000000000000;
    #10 assign a = 64'h51EFFFFFFFFFFFFF; assign b = 64'h6DFFFFFFFFFFFFFF;

    #10 $display("\n2**288 * 2**735:");
    #10 assign a = 64'h51F0000000000000; assign b = 64'h6DE0000000000000;
    #10 assign a = 64'h51FFFFFFFFFFFFFF; assign b = 64'h6DEFFFFFFFFFFFFF;

    #10 $display("\n2**289 * 2**734:");
    #10 assign a = 64'h5200000000000000; assign b = 64'h6DD0000000000000;
    #10 assign a = 64'h520FFFFFFFFFFFFF; assign b = 64'h6DDFFFFFFFFFFFFF;

    #10 $display("\n2**290 * 2**733:");
    #10 assign a = 64'h5210000000000000; assign b = 64'h6DC0000000000000;
    #10 assign a = 64'h521FFFFFFFFFFFFF; assign b = 64'h6DCFFFFFFFFFFFFF;

    #10 $display("\n2**291 * 2**732:");
    #10 assign a = 64'h5220000000000000; assign b = 64'h6DB0000000000000;
    #10 assign a = 64'h522FFFFFFFFFFFFF; assign b = 64'h6DBFFFFFFFFFFFFF;

    #10 $display("\n2**292 * 2**731:");
    #10 assign a = 64'h5230000000000000; assign b = 64'h6DA0000000000000;
    #10 assign a = 64'h523FFFFFFFFFFFFF; assign b = 64'h6DAFFFFFFFFFFFFF;

    #10 $display("\n2**293 * 2**730:");
    #10 assign a = 64'h5240000000000000; assign b = 64'h6D90000000000000;
    #10 assign a = 64'h524FFFFFFFFFFFFF; assign b = 64'h6D9FFFFFFFFFFFFF;

    #10 $display("\n2**294 * 2**729:");
    #10 assign a = 64'h5250000000000000; assign b = 64'h6D80000000000000;
    #10 assign a = 64'h525FFFFFFFFFFFFF; assign b = 64'h6D8FFFFFFFFFFFFF;

    #10 $display("\n2**295 * 2**728:");
    #10 assign a = 64'h5260000000000000; assign b = 64'h6D70000000000000;
    #10 assign a = 64'h526FFFFFFFFFFFFF; assign b = 64'h6D7FFFFFFFFFFFFF;

    #10 $display("\n2**296 * 2**727:");
    #10 assign a = 64'h5270000000000000; assign b = 64'h6D60000000000000;
    #10 assign a = 64'h527FFFFFFFFFFFFF; assign b = 64'h6D6FFFFFFFFFFFFF;

    #10 $display("\n2**297 * 2**726:");
    #10 assign a = 64'h5280000000000000; assign b = 64'h6D50000000000000;
    #10 assign a = 64'h528FFFFFFFFFFFFF; assign b = 64'h6D5FFFFFFFFFFFFF;

    #10 $display("\n2**298 * 2**725:");
    #10 assign a = 64'h5290000000000000; assign b = 64'h6D40000000000000;
    #10 assign a = 64'h529FFFFFFFFFFFFF; assign b = 64'h6D4FFFFFFFFFFFFF;

    #10 $display("\n2**299 * 2**724:");
    #10 assign a = 64'h52A0000000000000; assign b = 64'h6D30000000000000;
    #10 assign a = 64'h52AFFFFFFFFFFFFF; assign b = 64'h6D3FFFFFFFFFFFFF;

    #10 $display("\n2**300 * 2**723:");
    #10 assign a = 64'h52B0000000000000; assign b = 64'h6D20000000000000;
    #10 assign a = 64'h52BFFFFFFFFFFFFF; assign b = 64'h6D2FFFFFFFFFFFFF;

    #10 $display("\n2**301 * 2**722:");
    #10 assign a = 64'h52C0000000000000; assign b = 64'h6D10000000000000;
    #10 assign a = 64'h52CFFFFFFFFFFFFF; assign b = 64'h6D1FFFFFFFFFFFFF;

    #10 $display("\n2**302 * 2**721:");
    #10 assign a = 64'h52D0000000000000; assign b = 64'h6D00000000000000;
    #10 assign a = 64'h52DFFFFFFFFFFFFF; assign b = 64'h6D0FFFFFFFFFFFFF;

    #10 $display("\n2**303 * 2**720:");
    #10 assign a = 64'h52E0000000000000; assign b = 64'h6CF0000000000000;
    #10 assign a = 64'h52EFFFFFFFFFFFFF; assign b = 64'h6CFFFFFFFFFFFFFF;

    #10 $display("\n2**304 * 2**719:");
    #10 assign a = 64'h52F0000000000000; assign b = 64'h6CE0000000000000;
    #10 assign a = 64'h52FFFFFFFFFFFFFF; assign b = 64'h6CEFFFFFFFFFFFFF;

    #10 $display("\n2**305 * 2**718:");
    #10 assign a = 64'h5300000000000000; assign b = 64'h6CD0000000000000;
    #10 assign a = 64'h530FFFFFFFFFFFFF; assign b = 64'h6CDFFFFFFFFFFFFF;

    #10 $display("\n2**306 * 2**717:");
    #10 assign a = 64'h5310000000000000; assign b = 64'h6CC0000000000000;
    #10 assign a = 64'h531FFFFFFFFFFFFF; assign b = 64'h6CCFFFFFFFFFFFFF;

    #10 $display("\n2**307 * 2**716:");
    #10 assign a = 64'h5320000000000000; assign b = 64'h6CB0000000000000;
    #10 assign a = 64'h532FFFFFFFFFFFFF; assign b = 64'h6CBFFFFFFFFFFFFF;

    #10 $display("\n2**308 * 2**715:");
    #10 assign a = 64'h5330000000000000; assign b = 64'h6CA0000000000000;
    #10 assign a = 64'h533FFFFFFFFFFFFF; assign b = 64'h6CAFFFFFFFFFFFFF;

    #10 $display("\n2**309 * 2**714:");
    #10 assign a = 64'h5340000000000000; assign b = 64'h6C90000000000000;
    #10 assign a = 64'h534FFFFFFFFFFFFF; assign b = 64'h6C9FFFFFFFFFFFFF;

    #10 $display("\n2**310 * 2**713:");
    #10 assign a = 64'h5350000000000000; assign b = 64'h6C80000000000000;
    #10 assign a = 64'h535FFFFFFFFFFFFF; assign b = 64'h6C8FFFFFFFFFFFFF;

    #10 $display("\n2**311 * 2**712:");
    #10 assign a = 64'h5360000000000000; assign b = 64'h6C70000000000000;
    #10 assign a = 64'h536FFFFFFFFFFFFF; assign b = 64'h6C7FFFFFFFFFFFFF;

    #10 $display("\n2**312 * 2**711:");
    #10 assign a = 64'h5370000000000000; assign b = 64'h6C60000000000000;
    #10 assign a = 64'h537FFFFFFFFFFFFF; assign b = 64'h6C6FFFFFFFFFFFFF;

    #10 $display("\n2**313 * 2**710:");
    #10 assign a = 64'h5380000000000000; assign b = 64'h6C50000000000000;
    #10 assign a = 64'h538FFFFFFFFFFFFF; assign b = 64'h6C5FFFFFFFFFFFFF;

    #10 $display("\n2**314 * 2**709:");
    #10 assign a = 64'h5390000000000000; assign b = 64'h6C40000000000000;
    #10 assign a = 64'h539FFFFFFFFFFFFF; assign b = 64'h6C4FFFFFFFFFFFFF;

    #10 $display("\n2**315 * 2**708:");
    #10 assign a = 64'h53A0000000000000; assign b = 64'h6C30000000000000;
    #10 assign a = 64'h53AFFFFFFFFFFFFF; assign b = 64'h6C3FFFFFFFFFFFFF;

    #10 $display("\n2**316 * 2**707:");
    #10 assign a = 64'h53B0000000000000; assign b = 64'h6C20000000000000;
    #10 assign a = 64'h53BFFFFFFFFFFFFF; assign b = 64'h6C2FFFFFFFFFFFFF;

    #10 $display("\n2**317 * 2**706:");
    #10 assign a = 64'h53C0000000000000; assign b = 64'h6C10000000000000;
    #10 assign a = 64'h53CFFFFFFFFFFFFF; assign b = 64'h6C1FFFFFFFFFFFFF;

    #10 $display("\n2**318 * 2**705:");
    #10 assign a = 64'h53D0000000000000; assign b = 64'h6C00000000000000;
    #10 assign a = 64'h53DFFFFFFFFFFFFF; assign b = 64'h6C0FFFFFFFFFFFFF;

    #10 $display("\n2**319 * 2**704:");
    #10 assign a = 64'h53E0000000000000; assign b = 64'h6BF0000000000000;
    #10 assign a = 64'h53EFFFFFFFFFFFFF; assign b = 64'h6BFFFFFFFFFFFFFF;

    #10 $display("\n2**320 * 2**703:");
    #10 assign a = 64'h53F0000000000000; assign b = 64'h6BE0000000000000;
    #10 assign a = 64'h53FFFFFFFFFFFFFF; assign b = 64'h6BEFFFFFFFFFFFFF;

    #10 $display("\n2**321 * 2**702:");
    #10 assign a = 64'h5400000000000000; assign b = 64'h6BD0000000000000;
    #10 assign a = 64'h540FFFFFFFFFFFFF; assign b = 64'h6BDFFFFFFFFFFFFF;

    #10 $display("\n2**322 * 2**701:");
    #10 assign a = 64'h5410000000000000; assign b = 64'h6BC0000000000000;
    #10 assign a = 64'h541FFFFFFFFFFFFF; assign b = 64'h6BCFFFFFFFFFFFFF;

    #10 $display("\n2**323 * 2**700:");
    #10 assign a = 64'h5420000000000000; assign b = 64'h6BB0000000000000;
    #10 assign a = 64'h542FFFFFFFFFFFFF; assign b = 64'h6BBFFFFFFFFFFFFF;

    #10 $display("\n2**324 * 2**699:");
    #10 assign a = 64'h5430000000000000; assign b = 64'h6BA0000000000000;
    #10 assign a = 64'h543FFFFFFFFFFFFF; assign b = 64'h6BAFFFFFFFFFFFFF;

    #10 $display("\n2**325 * 2**698:");
    #10 assign a = 64'h5440000000000000; assign b = 64'h6B90000000000000;
    #10 assign a = 64'h544FFFFFFFFFFFFF; assign b = 64'h6B9FFFFFFFFFFFFF;

    #10 $display("\n2**326 * 2**697:");
    #10 assign a = 64'h5450000000000000; assign b = 64'h6B80000000000000;
    #10 assign a = 64'h545FFFFFFFFFFFFF; assign b = 64'h6B8FFFFFFFFFFFFF;

    #10 $display("\n2**327 * 2**696:");
    #10 assign a = 64'h5460000000000000; assign b = 64'h6B70000000000000;
    #10 assign a = 64'h546FFFFFFFFFFFFF; assign b = 64'h6B7FFFFFFFFFFFFF;

    #10 $display("\n2**328 * 2**695:");
    #10 assign a = 64'h5470000000000000; assign b = 64'h6B60000000000000;
    #10 assign a = 64'h547FFFFFFFFFFFFF; assign b = 64'h6B6FFFFFFFFFFFFF;

    #10 $display("\n2**329 * 2**694:");
    #10 assign a = 64'h5480000000000000; assign b = 64'h6B50000000000000;
    #10 assign a = 64'h548FFFFFFFFFFFFF; assign b = 64'h6B5FFFFFFFFFFFFF;

    #10 $display("\n2**330 * 2**693:");
    #10 assign a = 64'h5490000000000000; assign b = 64'h6B40000000000000;
    #10 assign a = 64'h549FFFFFFFFFFFFF; assign b = 64'h6B4FFFFFFFFFFFFF;

    #10 $display("\n2**331 * 2**692:");
    #10 assign a = 64'h54A0000000000000; assign b = 64'h6B30000000000000;
    #10 assign a = 64'h54AFFFFFFFFFFFFF; assign b = 64'h6B3FFFFFFFFFFFFF;

    #10 $display("\n2**332 * 2**691:");
    #10 assign a = 64'h54B0000000000000; assign b = 64'h6B20000000000000;
    #10 assign a = 64'h54BFFFFFFFFFFFFF; assign b = 64'h6B2FFFFFFFFFFFFF;

    #10 $display("\n2**333 * 2**690:");
    #10 assign a = 64'h54C0000000000000; assign b = 64'h6B10000000000000;
    #10 assign a = 64'h54CFFFFFFFFFFFFF; assign b = 64'h6B1FFFFFFFFFFFFF;

    #10 $display("\n2**334 * 2**689:");
    #10 assign a = 64'h54D0000000000000; assign b = 64'h6B00000000000000;
    #10 assign a = 64'h54DFFFFFFFFFFFFF; assign b = 64'h6B0FFFFFFFFFFFFF;

    #10 $display("\n2**335 * 2**688:");
    #10 assign a = 64'h54E0000000000000; assign b = 64'h6AF0000000000000;
    #10 assign a = 64'h54EFFFFFFFFFFFFF; assign b = 64'h6AFFFFFFFFFFFFFF;

    #10 $display("\n2**336 * 2**687:");
    #10 assign a = 64'h54F0000000000000; assign b = 64'h6AE0000000000000;
    #10 assign a = 64'h54FFFFFFFFFFFFFF; assign b = 64'h6AEFFFFFFFFFFFFF;

    #10 $display("\n2**337 * 2**686:");
    #10 assign a = 64'h5500000000000000; assign b = 64'h6AD0000000000000;
    #10 assign a = 64'h550FFFFFFFFFFFFF; assign b = 64'h6ADFFFFFFFFFFFFF;

    #10 $display("\n2**338 * 2**685:");
    #10 assign a = 64'h5510000000000000; assign b = 64'h6AC0000000000000;
    #10 assign a = 64'h551FFFFFFFFFFFFF; assign b = 64'h6ACFFFFFFFFFFFFF;

    #10 $display("\n2**339 * 2**684:");
    #10 assign a = 64'h5520000000000000; assign b = 64'h6AB0000000000000;
    #10 assign a = 64'h552FFFFFFFFFFFFF; assign b = 64'h6ABFFFFFFFFFFFFF;

    #10 $display("\n2**340 * 2**683:");
    #10 assign a = 64'h5530000000000000; assign b = 64'h6AA0000000000000;
    #10 assign a = 64'h553FFFFFFFFFFFFF; assign b = 64'h6AAFFFFFFFFFFFFF;

    #10 $display("\n2**341 * 2**682:");
    #10 assign a = 64'h5540000000000000; assign b = 64'h6A90000000000000;
    #10 assign a = 64'h554FFFFFFFFFFFFF; assign b = 64'h6A9FFFFFFFFFFFFF;

    #10 $display("\n2**342 * 2**681:");
    #10 assign a = 64'h5550000000000000; assign b = 64'h6A80000000000000;
    #10 assign a = 64'h555FFFFFFFFFFFFF; assign b = 64'h6A8FFFFFFFFFFFFF;

    #10 $display("\n2**343 * 2**680:");
    #10 assign a = 64'h5560000000000000; assign b = 64'h6A70000000000000;
    #10 assign a = 64'h556FFFFFFFFFFFFF; assign b = 64'h6A7FFFFFFFFFFFFF;

    #10 $display("\n2**344 * 2**679:");
    #10 assign a = 64'h5570000000000000; assign b = 64'h6A60000000000000;
    #10 assign a = 64'h557FFFFFFFFFFFFF; assign b = 64'h6A6FFFFFFFFFFFFF;

    #10 $display("\n2**345 * 2**678:");
    #10 assign a = 64'h5580000000000000; assign b = 64'h6A50000000000000;
    #10 assign a = 64'h558FFFFFFFFFFFFF; assign b = 64'h6A5FFFFFFFFFFFFF;

    #10 $display("\n2**346 * 2**677:");
    #10 assign a = 64'h5590000000000000; assign b = 64'h6A40000000000000;
    #10 assign a = 64'h559FFFFFFFFFFFFF; assign b = 64'h6A4FFFFFFFFFFFFF;

    #10 $display("\n2**347 * 2**676:");
    #10 assign a = 64'h55A0000000000000; assign b = 64'h6A30000000000000;
    #10 assign a = 64'h55AFFFFFFFFFFFFF; assign b = 64'h6A3FFFFFFFFFFFFF;

    #10 $display("\n2**348 * 2**675:");
    #10 assign a = 64'h55B0000000000000; assign b = 64'h6A20000000000000;
    #10 assign a = 64'h55BFFFFFFFFFFFFF; assign b = 64'h6A2FFFFFFFFFFFFF;

    #10 $display("\n2**349 * 2**674:");
    #10 assign a = 64'h55C0000000000000; assign b = 64'h6A10000000000000;
    #10 assign a = 64'h55CFFFFFFFFFFFFF; assign b = 64'h6A1FFFFFFFFFFFFF;

    #10 $display("\n2**350 * 2**673:");
    #10 assign a = 64'h55D0000000000000; assign b = 64'h6A00000000000000;
    #10 assign a = 64'h55DFFFFFFFFFFFFF; assign b = 64'h6A0FFFFFFFFFFFFF;

    #10 $display("\n2**351 * 2**672:");
    #10 assign a = 64'h55E0000000000000; assign b = 64'h69F0000000000000;
    #10 assign a = 64'h55EFFFFFFFFFFFFF; assign b = 64'h69FFFFFFFFFFFFFF;

    #10 $display("\n2**352 * 2**671:");
    #10 assign a = 64'h55F0000000000000; assign b = 64'h69E0000000000000;
    #10 assign a = 64'h55FFFFFFFFFFFFFF; assign b = 64'h69EFFFFFFFFFFFFF;

    #10 $display("\n2**353 * 2**670:");
    #10 assign a = 64'h5600000000000000; assign b = 64'h69D0000000000000;
    #10 assign a = 64'h560FFFFFFFFFFFFF; assign b = 64'h69DFFFFFFFFFFFFF;

    #10 $display("\n2**354 * 2**669:");
    #10 assign a = 64'h5610000000000000; assign b = 64'h69C0000000000000;
    #10 assign a = 64'h561FFFFFFFFFFFFF; assign b = 64'h69CFFFFFFFFFFFFF;

    #10 $display("\n2**355 * 2**668:");
    #10 assign a = 64'h5620000000000000; assign b = 64'h69B0000000000000;
    #10 assign a = 64'h562FFFFFFFFFFFFF; assign b = 64'h69BFFFFFFFFFFFFF;

    #10 $display("\n2**356 * 2**667:");
    #10 assign a = 64'h5630000000000000; assign b = 64'h69A0000000000000;
    #10 assign a = 64'h563FFFFFFFFFFFFF; assign b = 64'h69AFFFFFFFFFFFFF;

    #10 $display("\n2**357 * 2**666:");
    #10 assign a = 64'h5640000000000000; assign b = 64'h6990000000000000;
    #10 assign a = 64'h564FFFFFFFFFFFFF; assign b = 64'h699FFFFFFFFFFFFF;

    #10 $display("\n2**358 * 2**665:");
    #10 assign a = 64'h5650000000000000; assign b = 64'h6980000000000000;
    #10 assign a = 64'h565FFFFFFFFFFFFF; assign b = 64'h698FFFFFFFFFFFFF;

    #10 $display("\n2**359 * 2**664:");
    #10 assign a = 64'h5660000000000000; assign b = 64'h6970000000000000;
    #10 assign a = 64'h566FFFFFFFFFFFFF; assign b = 64'h697FFFFFFFFFFFFF;

    #10 $display("\n2**360 * 2**663:");
    #10 assign a = 64'h5670000000000000; assign b = 64'h6960000000000000;
    #10 assign a = 64'h567FFFFFFFFFFFFF; assign b = 64'h696FFFFFFFFFFFFF;

    #10 $display("\n2**361 * 2**662:");
    #10 assign a = 64'h5680000000000000; assign b = 64'h6950000000000000;
    #10 assign a = 64'h568FFFFFFFFFFFFF; assign b = 64'h695FFFFFFFFFFFFF;

    #10 $display("\n2**362 * 2**661:");
    #10 assign a = 64'h5690000000000000; assign b = 64'h6940000000000000;
    #10 assign a = 64'h569FFFFFFFFFFFFF; assign b = 64'h694FFFFFFFFFFFFF;

    #10 $display("\n2**363 * 2**660:");
    #10 assign a = 64'h56A0000000000000; assign b = 64'h6930000000000000;
    #10 assign a = 64'h56AFFFFFFFFFFFFF; assign b = 64'h693FFFFFFFFFFFFF;

    #10 $display("\n2**364 * 2**659:");
    #10 assign a = 64'h56B0000000000000; assign b = 64'h6920000000000000;
    #10 assign a = 64'h56BFFFFFFFFFFFFF; assign b = 64'h692FFFFFFFFFFFFF;

    #10 $display("\n2**365 * 2**658:");
    #10 assign a = 64'h56C0000000000000; assign b = 64'h6910000000000000;
    #10 assign a = 64'h56CFFFFFFFFFFFFF; assign b = 64'h691FFFFFFFFFFFFF;

    #10 $display("\n2**366 * 2**657:");
    #10 assign a = 64'h56D0000000000000; assign b = 64'h6900000000000000;
    #10 assign a = 64'h56DFFFFFFFFFFFFF; assign b = 64'h690FFFFFFFFFFFFF;

    #10 $display("\n2**367 * 2**656:");
    #10 assign a = 64'h56E0000000000000; assign b = 64'h68F0000000000000;
    #10 assign a = 64'h56EFFFFFFFFFFFFF; assign b = 64'h68FFFFFFFFFFFFFF;

    #10 $display("\n2**368 * 2**655:");
    #10 assign a = 64'h56F0000000000000; assign b = 64'h68E0000000000000;
    #10 assign a = 64'h56FFFFFFFFFFFFFF; assign b = 64'h68EFFFFFFFFFFFFF;

    #10 $display("\n2**369 * 2**654:");
    #10 assign a = 64'h5700000000000000; assign b = 64'h68D0000000000000;
    #10 assign a = 64'h570FFFFFFFFFFFFF; assign b = 64'h68DFFFFFFFFFFFFF;

    #10 $display("\n2**370 * 2**653:");
    #10 assign a = 64'h5710000000000000; assign b = 64'h68C0000000000000;
    #10 assign a = 64'h571FFFFFFFFFFFFF; assign b = 64'h68CFFFFFFFFFFFFF;

    #10 $display("\n2**371 * 2**652:");
    #10 assign a = 64'h5720000000000000; assign b = 64'h68B0000000000000;
    #10 assign a = 64'h572FFFFFFFFFFFFF; assign b = 64'h68BFFFFFFFFFFFFF;

    #10 $display("\n2**372 * 2**651:");
    #10 assign a = 64'h5730000000000000; assign b = 64'h68A0000000000000;
    #10 assign a = 64'h573FFFFFFFFFFFFF; assign b = 64'h68AFFFFFFFFFFFFF;

    #10 $display("\n2**373 * 2**650:");
    #10 assign a = 64'h5740000000000000; assign b = 64'h6890000000000000;
    #10 assign a = 64'h574FFFFFFFFFFFFF; assign b = 64'h689FFFFFFFFFFFFF;

    #10 $display("\n2**374 * 2**649:");
    #10 assign a = 64'h5750000000000000; assign b = 64'h6880000000000000;
    #10 assign a = 64'h575FFFFFFFFFFFFF; assign b = 64'h688FFFFFFFFFFFFF;

    #10 $display("\n2**375 * 2**648:");
    #10 assign a = 64'h5760000000000000; assign b = 64'h6870000000000000;
    #10 assign a = 64'h576FFFFFFFFFFFFF; assign b = 64'h687FFFFFFFFFFFFF;

    #10 $display("\n2**376 * 2**647:");
    #10 assign a = 64'h5770000000000000; assign b = 64'h6860000000000000;
    #10 assign a = 64'h577FFFFFFFFFFFFF; assign b = 64'h686FFFFFFFFFFFFF;

    #10 $display("\n2**377 * 2**646:");
    #10 assign a = 64'h5780000000000000; assign b = 64'h6850000000000000;
    #10 assign a = 64'h578FFFFFFFFFFFFF; assign b = 64'h685FFFFFFFFFFFFF;

    #10 $display("\n2**378 * 2**645:");
    #10 assign a = 64'h5790000000000000; assign b = 64'h6840000000000000;
    #10 assign a = 64'h579FFFFFFFFFFFFF; assign b = 64'h684FFFFFFFFFFFFF;

    #10 $display("\n2**379 * 2**644:");
    #10 assign a = 64'h57A0000000000000; assign b = 64'h6830000000000000;
    #10 assign a = 64'h57AFFFFFFFFFFFFF; assign b = 64'h683FFFFFFFFFFFFF;

    #10 $display("\n2**380 * 2**643:");
    #10 assign a = 64'h57B0000000000000; assign b = 64'h6820000000000000;
    #10 assign a = 64'h57BFFFFFFFFFFFFF; assign b = 64'h682FFFFFFFFFFFFF;

    #10 $display("\n2**381 * 2**642:");
    #10 assign a = 64'h57C0000000000000; assign b = 64'h6810000000000000;
    #10 assign a = 64'h57CFFFFFFFFFFFFF; assign b = 64'h681FFFFFFFFFFFFF;

    #10 $display("\n2**382 * 2**641:");
    #10 assign a = 64'h57D0000000000000; assign b = 64'h6800000000000000;
    #10 assign a = 64'h57DFFFFFFFFFFFFF; assign b = 64'h680FFFFFFFFFFFFF;

    #10 $display("\n2**383 * 2**640:");
    #10 assign a = 64'h57E0000000000000; assign b = 64'h67F0000000000000;
    #10 assign a = 64'h57EFFFFFFFFFFFFF; assign b = 64'h67FFFFFFFFFFFFFF;

    #10 $display("\n2**384 * 2**639:");
    #10 assign a = 64'h57F0000000000000; assign b = 64'h67E0000000000000;
    #10 assign a = 64'h57FFFFFFFFFFFFFF; assign b = 64'h67EFFFFFFFFFFFFF;

    #10 $display("\n2**385 * 2**638:");
    #10 assign a = 64'h5800000000000000; assign b = 64'h67D0000000000000;
    #10 assign a = 64'h580FFFFFFFFFFFFF; assign b = 64'h67DFFFFFFFFFFFFF;

    #10 $display("\n2**386 * 2**637:");
    #10 assign a = 64'h5810000000000000; assign b = 64'h67C0000000000000;
    #10 assign a = 64'h581FFFFFFFFFFFFF; assign b = 64'h67CFFFFFFFFFFFFF;

    #10 $display("\n2**387 * 2**636:");
    #10 assign a = 64'h5820000000000000; assign b = 64'h67B0000000000000;
    #10 assign a = 64'h582FFFFFFFFFFFFF; assign b = 64'h67BFFFFFFFFFFFFF;

    #10 $display("\n2**388 * 2**635:");
    #10 assign a = 64'h5830000000000000; assign b = 64'h67A0000000000000;
    #10 assign a = 64'h583FFFFFFFFFFFFF; assign b = 64'h67AFFFFFFFFFFFFF;

    #10 $display("\n2**389 * 2**634:");
    #10 assign a = 64'h5840000000000000; assign b = 64'h6790000000000000;
    #10 assign a = 64'h584FFFFFFFFFFFFF; assign b = 64'h679FFFFFFFFFFFFF;

    #10 $display("\n2**390 * 2**633:");
    #10 assign a = 64'h5850000000000000; assign b = 64'h6780000000000000;
    #10 assign a = 64'h585FFFFFFFFFFFFF; assign b = 64'h678FFFFFFFFFFFFF;

    #10 $display("\n2**391 * 2**632:");
    #10 assign a = 64'h5860000000000000; assign b = 64'h6770000000000000;
    #10 assign a = 64'h586FFFFFFFFFFFFF; assign b = 64'h677FFFFFFFFFFFFF;

    #10 $display("\n2**392 * 2**631:");
    #10 assign a = 64'h5870000000000000; assign b = 64'h6760000000000000;
    #10 assign a = 64'h587FFFFFFFFFFFFF; assign b = 64'h676FFFFFFFFFFFFF;

    #10 $display("\n2**393 * 2**630:");
    #10 assign a = 64'h5880000000000000; assign b = 64'h6750000000000000;
    #10 assign a = 64'h588FFFFFFFFFFFFF; assign b = 64'h675FFFFFFFFFFFFF;

    #10 $display("\n2**394 * 2**629:");
    #10 assign a = 64'h5890000000000000; assign b = 64'h6740000000000000;
    #10 assign a = 64'h589FFFFFFFFFFFFF; assign b = 64'h674FFFFFFFFFFFFF;

    #10 $display("\n2**395 * 2**628:");
    #10 assign a = 64'h58A0000000000000; assign b = 64'h6730000000000000;
    #10 assign a = 64'h58AFFFFFFFFFFFFF; assign b = 64'h673FFFFFFFFFFFFF;

    #10 $display("\n2**396 * 2**627:");
    #10 assign a = 64'h58B0000000000000; assign b = 64'h6720000000000000;
    #10 assign a = 64'h58BFFFFFFFFFFFFF; assign b = 64'h672FFFFFFFFFFFFF;

    #10 $display("\n2**397 * 2**626:");
    #10 assign a = 64'h58C0000000000000; assign b = 64'h6710000000000000;
    #10 assign a = 64'h58CFFFFFFFFFFFFF; assign b = 64'h671FFFFFFFFFFFFF;

    #10 $display("\n2**398 * 2**625:");
    #10 assign a = 64'h58D0000000000000; assign b = 64'h6700000000000000;
    #10 assign a = 64'h58DFFFFFFFFFFFFF; assign b = 64'h670FFFFFFFFFFFFF;

    #10 $display("\n2**399 * 2**624:");
    #10 assign a = 64'h58E0000000000000; assign b = 64'h66F0000000000000;
    #10 assign a = 64'h58EFFFFFFFFFFFFF; assign b = 64'h66FFFFFFFFFFFFFF;

    #10 $display("\n2**400 * 2**623:");
    #10 assign a = 64'h58F0000000000000; assign b = 64'h66E0000000000000;
    #10 assign a = 64'h58FFFFFFFFFFFFFF; assign b = 64'h66EFFFFFFFFFFFFF;

    #10 $display("\n2**401 * 2**622:");
    #10 assign a = 64'h5900000000000000; assign b = 64'h66D0000000000000;
    #10 assign a = 64'h590FFFFFFFFFFFFF; assign b = 64'h66DFFFFFFFFFFFFF;

    #10 $display("\n2**402 * 2**621:");
    #10 assign a = 64'h5910000000000000; assign b = 64'h66C0000000000000;
    #10 assign a = 64'h591FFFFFFFFFFFFF; assign b = 64'h66CFFFFFFFFFFFFF;

    #10 $display("\n2**403 * 2**620:");
    #10 assign a = 64'h5920000000000000; assign b = 64'h66B0000000000000;
    #10 assign a = 64'h592FFFFFFFFFFFFF; assign b = 64'h66BFFFFFFFFFFFFF;

    #10 $display("\n2**404 * 2**619:");
    #10 assign a = 64'h5930000000000000; assign b = 64'h66A0000000000000;
    #10 assign a = 64'h593FFFFFFFFFFFFF; assign b = 64'h66AFFFFFFFFFFFFF;

    #10 $display("\n2**405 * 2**618:");
    #10 assign a = 64'h5940000000000000; assign b = 64'h6690000000000000;
    #10 assign a = 64'h594FFFFFFFFFFFFF; assign b = 64'h669FFFFFFFFFFFFF;

    #10 $display("\n2**406 * 2**617:");
    #10 assign a = 64'h5950000000000000; assign b = 64'h6680000000000000;
    #10 assign a = 64'h595FFFFFFFFFFFFF; assign b = 64'h668FFFFFFFFFFFFF;

    #10 $display("\n2**407 * 2**616:");
    #10 assign a = 64'h5960000000000000; assign b = 64'h6670000000000000;
    #10 assign a = 64'h596FFFFFFFFFFFFF; assign b = 64'h667FFFFFFFFFFFFF;

    #10 $display("\n2**408 * 2**615:");
    #10 assign a = 64'h5970000000000000; assign b = 64'h6660000000000000;
    #10 assign a = 64'h597FFFFFFFFFFFFF; assign b = 64'h666FFFFFFFFFFFFF;

    #10 $display("\n2**409 * 2**614:");
    #10 assign a = 64'h5980000000000000; assign b = 64'h6650000000000000;
    #10 assign a = 64'h598FFFFFFFFFFFFF; assign b = 64'h665FFFFFFFFFFFFF;

    #10 $display("\n2**410 * 2**613:");
    #10 assign a = 64'h5990000000000000; assign b = 64'h6640000000000000;
    #10 assign a = 64'h599FFFFFFFFFFFFF; assign b = 64'h664FFFFFFFFFFFFF;

    #10 $display("\n2**411 * 2**612:");
    #10 assign a = 64'h59A0000000000000; assign b = 64'h6630000000000000;
    #10 assign a = 64'h59AFFFFFFFFFFFFF; assign b = 64'h663FFFFFFFFFFFFF;

    #10 $display("\n2**412 * 2**611:");
    #10 assign a = 64'h59B0000000000000; assign b = 64'h6620000000000000;
    #10 assign a = 64'h59BFFFFFFFFFFFFF; assign b = 64'h662FFFFFFFFFFFFF;

    #10 $display("\n2**413 * 2**610:");
    #10 assign a = 64'h59C0000000000000; assign b = 64'h6610000000000000;
    #10 assign a = 64'h59CFFFFFFFFFFFFF; assign b = 64'h661FFFFFFFFFFFFF;

    #10 $display("\n2**414 * 2**609:");
    #10 assign a = 64'h59D0000000000000; assign b = 64'h6600000000000000;
    #10 assign a = 64'h59DFFFFFFFFFFFFF; assign b = 64'h660FFFFFFFFFFFFF;

    #10 $display("\n2**415 * 2**608:");
    #10 assign a = 64'h59E0000000000000; assign b = 64'h65F0000000000000;
    #10 assign a = 64'h59EFFFFFFFFFFFFF; assign b = 64'h65FFFFFFFFFFFFFF;

    #10 $display("\n2**416 * 2**607:");
    #10 assign a = 64'h59F0000000000000; assign b = 64'h65E0000000000000;
    #10 assign a = 64'h59FFFFFFFFFFFFFF; assign b = 64'h65EFFFFFFFFFFFFF;

    #10 $display("\n2**417 * 2**606:");
    #10 assign a = 64'h5A00000000000000; assign b = 64'h65D0000000000000;
    #10 assign a = 64'h5A0FFFFFFFFFFFFF; assign b = 64'h65DFFFFFFFFFFFFF;

    #10 $display("\n2**418 * 2**605:");
    #10 assign a = 64'h5A10000000000000; assign b = 64'h65C0000000000000;
    #10 assign a = 64'h5A1FFFFFFFFFFFFF; assign b = 64'h65CFFFFFFFFFFFFF;

    #10 $display("\n2**419 * 2**604:");
    #10 assign a = 64'h5A20000000000000; assign b = 64'h65B0000000000000;
    #10 assign a = 64'h5A2FFFFFFFFFFFFF; assign b = 64'h65BFFFFFFFFFFFFF;

    #10 $display("\n2**420 * 2**603:");
    #10 assign a = 64'h5A30000000000000; assign b = 64'h65A0000000000000;
    #10 assign a = 64'h5A3FFFFFFFFFFFFF; assign b = 64'h65AFFFFFFFFFFFFF;

    #10 $display("\n2**421 * 2**602:");
    #10 assign a = 64'h5A40000000000000; assign b = 64'h6590000000000000;
    #10 assign a = 64'h5A4FFFFFFFFFFFFF; assign b = 64'h659FFFFFFFFFFFFF;

    #10 $display("\n2**422 * 2**601:");
    #10 assign a = 64'h5A50000000000000; assign b = 64'h6580000000000000;
    #10 assign a = 64'h5A5FFFFFFFFFFFFF; assign b = 64'h658FFFFFFFFFFFFF;

    #10 $display("\n2**423 * 2**600:");
    #10 assign a = 64'h5A60000000000000; assign b = 64'h6570000000000000;
    #10 assign a = 64'h5A6FFFFFFFFFFFFF; assign b = 64'h657FFFFFFFFFFFFF;

    #10 $display("\n2**424 * 2**599:");
    #10 assign a = 64'h5A70000000000000; assign b = 64'h6560000000000000;
    #10 assign a = 64'h5A7FFFFFFFFFFFFF; assign b = 64'h656FFFFFFFFFFFFF;

    #10 $display("\n2**425 * 2**598:");
    #10 assign a = 64'h5A80000000000000; assign b = 64'h6550000000000000;
    #10 assign a = 64'h5A8FFFFFFFFFFFFF; assign b = 64'h655FFFFFFFFFFFFF;

    #10 $display("\n2**426 * 2**597:");
    #10 assign a = 64'h5A90000000000000; assign b = 64'h6540000000000000;
    #10 assign a = 64'h5A9FFFFFFFFFFFFF; assign b = 64'h654FFFFFFFFFFFFF;

    #10 $display("\n2**427 * 2**596:");
    #10 assign a = 64'h5AA0000000000000; assign b = 64'h6530000000000000;
    #10 assign a = 64'h5AAFFFFFFFFFFFFF; assign b = 64'h653FFFFFFFFFFFFF;

    #10 $display("\n2**428 * 2**595:");
    #10 assign a = 64'h5AB0000000000000; assign b = 64'h6520000000000000;
    #10 assign a = 64'h5ABFFFFFFFFFFFFF; assign b = 64'h652FFFFFFFFFFFFF;

    #10 $display("\n2**429 * 2**594:");
    #10 assign a = 64'h5AC0000000000000; assign b = 64'h6510000000000000;
    #10 assign a = 64'h5ACFFFFFFFFFFFFF; assign b = 64'h651FFFFFFFFFFFFF;

    #10 $display("\n2**430 * 2**593:");
    #10 assign a = 64'h5AD0000000000000; assign b = 64'h6500000000000000;
    #10 assign a = 64'h5ADFFFFFFFFFFFFF; assign b = 64'h650FFFFFFFFFFFFF;

    #10 $display("\n2**431 * 2**592:");
    #10 assign a = 64'h5AE0000000000000; assign b = 64'h64F0000000000000;
    #10 assign a = 64'h5AEFFFFFFFFFFFFF; assign b = 64'h64FFFFFFFFFFFFFF;

    #10 $display("\n2**432 * 2**591:");
    #10 assign a = 64'h5AF0000000000000; assign b = 64'h64E0000000000000;
    #10 assign a = 64'h5AFFFFFFFFFFFFFF; assign b = 64'h64EFFFFFFFFFFFFF;

    #10 $display("\n2**433 * 2**590:");
    #10 assign a = 64'h5B00000000000000; assign b = 64'h64D0000000000000;
    #10 assign a = 64'h5B0FFFFFFFFFFFFF; assign b = 64'h64DFFFFFFFFFFFFF;

    #10 $display("\n2**434 * 2**589:");
    #10 assign a = 64'h5B10000000000000; assign b = 64'h64C0000000000000;
    #10 assign a = 64'h5B1FFFFFFFFFFFFF; assign b = 64'h64CFFFFFFFFFFFFF;

    #10 $display("\n2**435 * 2**588:");
    #10 assign a = 64'h5B20000000000000; assign b = 64'h64B0000000000000;
    #10 assign a = 64'h5B2FFFFFFFFFFFFF; assign b = 64'h64BFFFFFFFFFFFFF;

    #10 $display("\n2**436 * 2**587:");
    #10 assign a = 64'h5B30000000000000; assign b = 64'h64A0000000000000;
    #10 assign a = 64'h5B3FFFFFFFFFFFFF; assign b = 64'h64AFFFFFFFFFFFFF;

    #10 $display("\n2**437 * 2**586:");
    #10 assign a = 64'h5B40000000000000; assign b = 64'h6490000000000000;
    #10 assign a = 64'h5B4FFFFFFFFFFFFF; assign b = 64'h649FFFFFFFFFFFFF;

    #10 $display("\n2**438 * 2**585:");
    #10 assign a = 64'h5B50000000000000; assign b = 64'h6480000000000000;
    #10 assign a = 64'h5B5FFFFFFFFFFFFF; assign b = 64'h648FFFFFFFFFFFFF;

    #10 $display("\n2**439 * 2**584:");
    #10 assign a = 64'h5B60000000000000; assign b = 64'h6470000000000000;
    #10 assign a = 64'h5B6FFFFFFFFFFFFF; assign b = 64'h647FFFFFFFFFFFFF;

    #10 $display("\n2**440 * 2**583:");
    #10 assign a = 64'h5B70000000000000; assign b = 64'h6460000000000000;
    #10 assign a = 64'h5B7FFFFFFFFFFFFF; assign b = 64'h646FFFFFFFFFFFFF;

    #10 $display("\n2**441 * 2**582:");
    #10 assign a = 64'h5B80000000000000; assign b = 64'h6450000000000000;
    #10 assign a = 64'h5B8FFFFFFFFFFFFF; assign b = 64'h645FFFFFFFFFFFFF;

    #10 $display("\n2**442 * 2**581:");
    #10 assign a = 64'h5B90000000000000; assign b = 64'h6440000000000000;
    #10 assign a = 64'h5B9FFFFFFFFFFFFF; assign b = 64'h644FFFFFFFFFFFFF;

    #10 $display("\n2**443 * 2**580:");
    #10 assign a = 64'h5BA0000000000000; assign b = 64'h6430000000000000;
    #10 assign a = 64'h5BAFFFFFFFFFFFFF; assign b = 64'h643FFFFFFFFFFFFF;

    #10 $display("\n2**444 * 2**579:");
    #10 assign a = 64'h5BB0000000000000; assign b = 64'h6420000000000000;
    #10 assign a = 64'h5BBFFFFFFFFFFFFF; assign b = 64'h642FFFFFFFFFFFFF;

    #10 $display("\n2**445 * 2**578:");
    #10 assign a = 64'h5BC0000000000000; assign b = 64'h6410000000000000;
    #10 assign a = 64'h5BCFFFFFFFFFFFFF; assign b = 64'h641FFFFFFFFFFFFF;

    #10 $display("\n2**446 * 2**577:");
    #10 assign a = 64'h5BD0000000000000; assign b = 64'h6400000000000000;
    #10 assign a = 64'h5BDFFFFFFFFFFFFF; assign b = 64'h640FFFFFFFFFFFFF;

    #10 $display("\n2**447 * 2**576:");
    #10 assign a = 64'h5BE0000000000000; assign b = 64'h63F0000000000000;
    #10 assign a = 64'h5BEFFFFFFFFFFFFF; assign b = 64'h63FFFFFFFFFFFFFF;

    #10 $display("\n2**448 * 2**575:");
    #10 assign a = 64'h5BF0000000000000; assign b = 64'h63E0000000000000;
    #10 assign a = 64'h5BFFFFFFFFFFFFFF; assign b = 64'h63EFFFFFFFFFFFFF;

    #10 $display("\n2**449 * 2**574:");
    #10 assign a = 64'h5C00000000000000; assign b = 64'h63D0000000000000;
    #10 assign a = 64'h5C0FFFFFFFFFFFFF; assign b = 64'h63DFFFFFFFFFFFFF;

    #10 $display("\n2**450 * 2**573:");
    #10 assign a = 64'h5C10000000000000; assign b = 64'h63C0000000000000;
    #10 assign a = 64'h5C1FFFFFFFFFFFFF; assign b = 64'h63CFFFFFFFFFFFFF;

    #10 $display("\n2**451 * 2**572:");
    #10 assign a = 64'h5C20000000000000; assign b = 64'h63B0000000000000;
    #10 assign a = 64'h5C2FFFFFFFFFFFFF; assign b = 64'h63BFFFFFFFFFFFFF;

    #10 $display("\n2**452 * 2**571:");
    #10 assign a = 64'h5C30000000000000; assign b = 64'h63A0000000000000;
    #10 assign a = 64'h5C3FFFFFFFFFFFFF; assign b = 64'h63AFFFFFFFFFFFFF;

    #10 $display("\n2**453 * 2**570:");
    #10 assign a = 64'h5C40000000000000; assign b = 64'h6390000000000000;
    #10 assign a = 64'h5C4FFFFFFFFFFFFF; assign b = 64'h639FFFFFFFFFFFFF;

    #10 $display("\n2**454 * 2**569:");
    #10 assign a = 64'h5C50000000000000; assign b = 64'h6380000000000000;
    #10 assign a = 64'h5C5FFFFFFFFFFFFF; assign b = 64'h638FFFFFFFFFFFFF;

    #10 $display("\n2**455 * 2**568:");
    #10 assign a = 64'h5C60000000000000; assign b = 64'h6370000000000000;
    #10 assign a = 64'h5C6FFFFFFFFFFFFF; assign b = 64'h637FFFFFFFFFFFFF;

    #10 $display("\n2**456 * 2**567:");
    #10 assign a = 64'h5C70000000000000; assign b = 64'h6360000000000000;
    #10 assign a = 64'h5C7FFFFFFFFFFFFF; assign b = 64'h636FFFFFFFFFFFFF;

    #10 $display("\n2**457 * 2**566:");
    #10 assign a = 64'h5C80000000000000; assign b = 64'h6350000000000000;
    #10 assign a = 64'h5C8FFFFFFFFFFFFF; assign b = 64'h635FFFFFFFFFFFFF;

    #10 $display("\n2**458 * 2**565:");
    #10 assign a = 64'h5C90000000000000; assign b = 64'h6340000000000000;
    #10 assign a = 64'h5C9FFFFFFFFFFFFF; assign b = 64'h634FFFFFFFFFFFFF;

    #10 $display("\n2**459 * 2**564:");
    #10 assign a = 64'h5CA0000000000000; assign b = 64'h6330000000000000;
    #10 assign a = 64'h5CAFFFFFFFFFFFFF; assign b = 64'h633FFFFFFFFFFFFF;

    #10 $display("\n2**460 * 2**563:");
    #10 assign a = 64'h5CB0000000000000; assign b = 64'h6320000000000000;
    #10 assign a = 64'h5CBFFFFFFFFFFFFF; assign b = 64'h632FFFFFFFFFFFFF;

    #10 $display("\n2**461 * 2**562:");
    #10 assign a = 64'h5CC0000000000000; assign b = 64'h6310000000000000;
    #10 assign a = 64'h5CCFFFFFFFFFFFFF; assign b = 64'h631FFFFFFFFFFFFF;

    #10 $display("\n2**462 * 2**561:");
    #10 assign a = 64'h5CD0000000000000; assign b = 64'h6300000000000000;
    #10 assign a = 64'h5CDFFFFFFFFFFFFF; assign b = 64'h630FFFFFFFFFFFFF;

    #10 $display("\n2**463 * 2**560:");
    #10 assign a = 64'h5CE0000000000000; assign b = 64'h62F0000000000000;
    #10 assign a = 64'h5CEFFFFFFFFFFFFF; assign b = 64'h62FFFFFFFFFFFFFF;

    #10 $display("\n2**464 * 2**559:");
    #10 assign a = 64'h5CF0000000000000; assign b = 64'h62E0000000000000;
    #10 assign a = 64'h5CFFFFFFFFFFFFFF; assign b = 64'h62EFFFFFFFFFFFFF;

    #10 $display("\n2**465 * 2**558:");
    #10 assign a = 64'h5D00000000000000; assign b = 64'h62D0000000000000;
    #10 assign a = 64'h5D0FFFFFFFFFFFFF; assign b = 64'h62DFFFFFFFFFFFFF;

    #10 $display("\n2**466 * 2**557:");
    #10 assign a = 64'h5D10000000000000; assign b = 64'h62C0000000000000;
    #10 assign a = 64'h5D1FFFFFFFFFFFFF; assign b = 64'h62CFFFFFFFFFFFFF;

    #10 $display("\n2**467 * 2**556:");
    #10 assign a = 64'h5D20000000000000; assign b = 64'h62B0000000000000;
    #10 assign a = 64'h5D2FFFFFFFFFFFFF; assign b = 64'h62BFFFFFFFFFFFFF;

    #10 $display("\n2**468 * 2**555:");
    #10 assign a = 64'h5D30000000000000; assign b = 64'h62A0000000000000;
    #10 assign a = 64'h5D3FFFFFFFFFFFFF; assign b = 64'h62AFFFFFFFFFFFFF;

    #10 $display("\n2**469 * 2**554:");
    #10 assign a = 64'h5D40000000000000; assign b = 64'h6290000000000000;
    #10 assign a = 64'h5D4FFFFFFFFFFFFF; assign b = 64'h629FFFFFFFFFFFFF;

    #10 $display("\n2**470 * 2**553:");
    #10 assign a = 64'h5D50000000000000; assign b = 64'h6280000000000000;
    #10 assign a = 64'h5D5FFFFFFFFFFFFF; assign b = 64'h628FFFFFFFFFFFFF;

    #10 $display("\n2**471 * 2**552:");
    #10 assign a = 64'h5D60000000000000; assign b = 64'h6270000000000000;
    #10 assign a = 64'h5D6FFFFFFFFFFFFF; assign b = 64'h627FFFFFFFFFFFFF;

    #10 $display("\n2**472 * 2**551:");
    #10 assign a = 64'h5D70000000000000; assign b = 64'h6260000000000000;
    #10 assign a = 64'h5D7FFFFFFFFFFFFF; assign b = 64'h626FFFFFFFFFFFFF;

    #10 $display("\n2**473 * 2**550:");
    #10 assign a = 64'h5D80000000000000; assign b = 64'h6250000000000000;
    #10 assign a = 64'h5D8FFFFFFFFFFFFF; assign b = 64'h625FFFFFFFFFFFFF;

    #10 $display("\n2**474 * 2**549:");
    #10 assign a = 64'h5D90000000000000; assign b = 64'h6240000000000000;
    #10 assign a = 64'h5D9FFFFFFFFFFFFF; assign b = 64'h624FFFFFFFFFFFFF;

    #10 $display("\n2**475 * 2**548:");
    #10 assign a = 64'h5DA0000000000000; assign b = 64'h6230000000000000;
    #10 assign a = 64'h5DAFFFFFFFFFFFFF; assign b = 64'h623FFFFFFFFFFFFF;

    #10 $display("\n2**476 * 2**547:");
    #10 assign a = 64'h5DB0000000000000; assign b = 64'h6220000000000000;
    #10 assign a = 64'h5DBFFFFFFFFFFFFF; assign b = 64'h622FFFFFFFFFFFFF;

    #10 $display("\n2**477 * 2**546:");
    #10 assign a = 64'h5DC0000000000000; assign b = 64'h6210000000000000;
    #10 assign a = 64'h5DCFFFFFFFFFFFFF; assign b = 64'h621FFFFFFFFFFFFF;

    #10 $display("\n2**478 * 2**545:");
    #10 assign a = 64'h5DD0000000000000; assign b = 64'h6200000000000000;
    #10 assign a = 64'h5DDFFFFFFFFFFFFF; assign b = 64'h620FFFFFFFFFFFFF;

    #10 $display("\n2**479 * 2**544:");
    #10 assign a = 64'h5DE0000000000000; assign b = 64'h61F0000000000000;
    #10 assign a = 64'h5DEFFFFFFFFFFFFF; assign b = 64'h61FFFFFFFFFFFFFF;

    #10 $display("\n2**480 * 2**543:");
    #10 assign a = 64'h5DF0000000000000; assign b = 64'h61E0000000000000;
    #10 assign a = 64'h5DFFFFFFFFFFFFFF; assign b = 64'h61EFFFFFFFFFFFFF;

    #10 $display("\n2**481 * 2**542:");
    #10 assign a = 64'h5E00000000000000; assign b = 64'h61D0000000000000;
    #10 assign a = 64'h5E0FFFFFFFFFFFFF; assign b = 64'h61DFFFFFFFFFFFFF;

    #10 $display("\n2**482 * 2**541:");
    #10 assign a = 64'h5E10000000000000; assign b = 64'h61C0000000000000;
    #10 assign a = 64'h5E1FFFFFFFFFFFFF; assign b = 64'h61CFFFFFFFFFFFFF;

    #10 $display("\n2**483 * 2**540:");
    #10 assign a = 64'h5E20000000000000; assign b = 64'h61B0000000000000;
    #10 assign a = 64'h5E2FFFFFFFFFFFFF; assign b = 64'h61BFFFFFFFFFFFFF;

    #10 $display("\n2**484 * 2**539:");
    #10 assign a = 64'h5E30000000000000; assign b = 64'h61A0000000000000;
    #10 assign a = 64'h5E3FFFFFFFFFFFFF; assign b = 64'h61AFFFFFFFFFFFFF;

    #10 $display("\n2**485 * 2**538:");
    #10 assign a = 64'h5E40000000000000; assign b = 64'h6190000000000000;
    #10 assign a = 64'h5E4FFFFFFFFFFFFF; assign b = 64'h619FFFFFFFFFFFFF;

    #10 $display("\n2**486 * 2**537:");
    #10 assign a = 64'h5E50000000000000; assign b = 64'h6180000000000000;
    #10 assign a = 64'h5E5FFFFFFFFFFFFF; assign b = 64'h618FFFFFFFFFFFFF;

    #10 $display("\n2**487 * 2**536:");
    #10 assign a = 64'h5E60000000000000; assign b = 64'h6170000000000000;
    #10 assign a = 64'h5E6FFFFFFFFFFFFF; assign b = 64'h617FFFFFFFFFFFFF;

    #10 $display("\n2**488 * 2**535:");
    #10 assign a = 64'h5E70000000000000; assign b = 64'h6160000000000000;
    #10 assign a = 64'h5E7FFFFFFFFFFFFF; assign b = 64'h616FFFFFFFFFFFFF;

    #10 $display("\n2**489 * 2**534:");
    #10 assign a = 64'h5E80000000000000; assign b = 64'h6150000000000000;
    #10 assign a = 64'h5E8FFFFFFFFFFFFF; assign b = 64'h615FFFFFFFFFFFFF;

    #10 $display("\n2**490 * 2**533:");
    #10 assign a = 64'h5E90000000000000; assign b = 64'h6140000000000000;
    #10 assign a = 64'h5E9FFFFFFFFFFFFF; assign b = 64'h614FFFFFFFFFFFFF;

    #10 $display("\n2**491 * 2**532:");
    #10 assign a = 64'h5EA0000000000000; assign b = 64'h6130000000000000;
    #10 assign a = 64'h5EAFFFFFFFFFFFFF; assign b = 64'h613FFFFFFFFFFFFF;

    #10 $display("\n2**492 * 2**531:");
    #10 assign a = 64'h5EB0000000000000; assign b = 64'h6120000000000000;
    #10 assign a = 64'h5EBFFFFFFFFFFFFF; assign b = 64'h612FFFFFFFFFFFFF;

    #10 $display("\n2**493 * 2**530:");
    #10 assign a = 64'h5EC0000000000000; assign b = 64'h6110000000000000;
    #10 assign a = 64'h5ECFFFFFFFFFFFFF; assign b = 64'h611FFFFFFFFFFFFF;

    #10 $display("\n2**494 * 2**529:");
    #10 assign a = 64'h5ED0000000000000; assign b = 64'h6100000000000000;
    #10 assign a = 64'h5EDFFFFFFFFFFFFF; assign b = 64'h610FFFFFFFFFFFFF;

    #10 $display("\n2**495 * 2**528:");
    #10 assign a = 64'h5EE0000000000000; assign b = 64'h60F0000000000000;
    #10 assign a = 64'h5EEFFFFFFFFFFFFF; assign b = 64'h60FFFFFFFFFFFFFF;

    #10 $display("\n2**496 * 2**527:");
    #10 assign a = 64'h5EF0000000000000; assign b = 64'h60E0000000000000;
    #10 assign a = 64'h5EFFFFFFFFFFFFFF; assign b = 64'h60EFFFFFFFFFFFFF;

    #10 $display("\n2**497 * 2**526:");
    #10 assign a = 64'h5F00000000000000; assign b = 64'h60D0000000000000;
    #10 assign a = 64'h5F0FFFFFFFFFFFFF; assign b = 64'h60DFFFFFFFFFFFFF;

    #10 $display("\n2**498 * 2**525:");
    #10 assign a = 64'h5F10000000000000; assign b = 64'h60C0000000000000;
    #10 assign a = 64'h5F1FFFFFFFFFFFFF; assign b = 64'h60CFFFFFFFFFFFFF;

    #10 $display("\n2**499 * 2**524:");
    #10 assign a = 64'h5F20000000000000; assign b = 64'h60B0000000000000;
    #10 assign a = 64'h5F2FFFFFFFFFFFFF; assign b = 64'h60BFFFFFFFFFFFFF;

    #10 $display("\n2**500 * 2**523:");
    #10 assign a = 64'h5F30000000000000; assign b = 64'h60A0000000000000;
    #10 assign a = 64'h5F3FFFFFFFFFFFFF; assign b = 64'h60AFFFFFFFFFFFFF;

    #10 $display("\n2**501 * 2**522:");
    #10 assign a = 64'h5F40000000000000; assign b = 64'h6090000000000000;
    #10 assign a = 64'h5F4FFFFFFFFFFFFF; assign b = 64'h609FFFFFFFFFFFFF;

    #10 $display("\n2**502 * 2**521:");
    #10 assign a = 64'h5F50000000000000; assign b = 64'h6080000000000000;
    #10 assign a = 64'h5F5FFFFFFFFFFFFF; assign b = 64'h608FFFFFFFFFFFFF;

    #10 $display("\n2**503 * 2**520:");
    #10 assign a = 64'h5F60000000000000; assign b = 64'h6070000000000000;
    #10 assign a = 64'h5F6FFFFFFFFFFFFF; assign b = 64'h607FFFFFFFFFFFFF;

    #10 $display("\n2**504 * 2**519:");
    #10 assign a = 64'h5F70000000000000; assign b = 64'h6060000000000000;
    #10 assign a = 64'h5F7FFFFFFFFFFFFF; assign b = 64'h606FFFFFFFFFFFFF;

    #10 $display("\n2**505 * 2**518:");
    #10 assign a = 64'h5F80000000000000; assign b = 64'h6050000000000000;
    #10 assign a = 64'h5F8FFFFFFFFFFFFF; assign b = 64'h605FFFFFFFFFFFFF;

    #10 $display("\n2**506 * 2**517:");
    #10 assign a = 64'h5F90000000000000; assign b = 64'h6040000000000000;
    #10 assign a = 64'h5F9FFFFFFFFFFFFF; assign b = 64'h604FFFFFFFFFFFFF;

    #10 $display("\n2**507 * 2**516:");
    #10 assign a = 64'h5FA0000000000000; assign b = 64'h6030000000000000;
    #10 assign a = 64'h5FAFFFFFFFFFFFFF; assign b = 64'h603FFFFFFFFFFFFF;

    #10 $display("\n2**508 * 2**515:");
    #10 assign a = 64'h5FB0000000000000; assign b = 64'h6020000000000000;
    #10 assign a = 64'h5FBFFFFFFFFFFFFF; assign b = 64'h602FFFFFFFFFFFFF;

    #10 $display("\n2**509 * 2**514:");
    #10 assign a = 64'h5FC0000000000000; assign b = 64'h6010000000000000;
    #10 assign a = 64'h5FCFFFFFFFFFFFFF; assign b = 64'h601FFFFFFFFFFFFF;

    #10 $display("\n2**510 * 2**513:");
    #10 assign a = 64'h5FD0000000000000; assign b = 64'h6000000000000000;
    #10 assign a = 64'h5FDFFFFFFFFFFFFF; assign b = 64'h600FFFFFFFFFFFFF;

    #10 $display("\n2**511 * 2**512:");
    #10 assign a = 64'h5FE0000000000000; assign b = 64'h5FF0000000000000;
    #10 assign a = 64'h5FEFFFFFFFFFFFFF; assign b = 64'h5FFFFFFFFFFFFFFF;

    #10 $display("\n2**512 * 2**511:");
    #10 assign a = 64'h5FF0000000000000; assign b = 64'h5FE0000000000000;
    #10 assign a = 64'h5FFFFFFFFFFFFFFF; assign b = 64'h5FEFFFFFFFFFFFFF;

    #10 $display("\n2**513 * 2**510:");
    #10 assign a = 64'h6000000000000000; assign b = 64'h5FD0000000000000;
    #10 assign a = 64'h600FFFFFFFFFFFFF; assign b = 64'h5FDFFFFFFFFFFFFF;

    #10 $display("\n2**514 * 2**509:");
    #10 assign a = 64'h6010000000000000; assign b = 64'h5FC0000000000000;
    #10 assign a = 64'h601FFFFFFFFFFFFF; assign b = 64'h5FCFFFFFFFFFFFFF;

    #10 $display("\n2**515 * 2**508:");
    #10 assign a = 64'h6020000000000000; assign b = 64'h5FB0000000000000;
    #10 assign a = 64'h602FFFFFFFFFFFFF; assign b = 64'h5FBFFFFFFFFFFFFF;

    #10 $display("\n2**516 * 2**507:");
    #10 assign a = 64'h6030000000000000; assign b = 64'h5FA0000000000000;
    #10 assign a = 64'h603FFFFFFFFFFFFF; assign b = 64'h5FAFFFFFFFFFFFFF;

    #10 $display("\n2**517 * 2**506:");
    #10 assign a = 64'h6040000000000000; assign b = 64'h5F90000000000000;
    #10 assign a = 64'h604FFFFFFFFFFFFF; assign b = 64'h5F9FFFFFFFFFFFFF;

    #10 $display("\n2**518 * 2**505:");
    #10 assign a = 64'h6050000000000000; assign b = 64'h5F80000000000000;
    #10 assign a = 64'h605FFFFFFFFFFFFF; assign b = 64'h5F8FFFFFFFFFFFFF;

    #10 $display("\n2**519 * 2**504:");
    #10 assign a = 64'h6060000000000000; assign b = 64'h5F70000000000000;
    #10 assign a = 64'h606FFFFFFFFFFFFF; assign b = 64'h5F7FFFFFFFFFFFFF;

    #10 $display("\n2**520 * 2**503:");
    #10 assign a = 64'h6070000000000000; assign b = 64'h5F60000000000000;
    #10 assign a = 64'h607FFFFFFFFFFFFF; assign b = 64'h5F6FFFFFFFFFFFFF;

    #10 $display("\n2**521 * 2**502:");
    #10 assign a = 64'h6080000000000000; assign b = 64'h5F50000000000000;
    #10 assign a = 64'h608FFFFFFFFFFFFF; assign b = 64'h5F5FFFFFFFFFFFFF;

    #10 $display("\n2**522 * 2**501:");
    #10 assign a = 64'h6090000000000000; assign b = 64'h5F40000000000000;
    #10 assign a = 64'h609FFFFFFFFFFFFF; assign b = 64'h5F4FFFFFFFFFFFFF;

    #10 $display("\n2**523 * 2**500:");
    #10 assign a = 64'h60A0000000000000; assign b = 64'h5F30000000000000;
    #10 assign a = 64'h60AFFFFFFFFFFFFF; assign b = 64'h5F3FFFFFFFFFFFFF;

    #10 $display("\n2**524 * 2**499:");
    #10 assign a = 64'h60B0000000000000; assign b = 64'h5F20000000000000;
    #10 assign a = 64'h60BFFFFFFFFFFFFF; assign b = 64'h5F2FFFFFFFFFFFFF;

    #10 $display("\n2**525 * 2**498:");
    #10 assign a = 64'h60C0000000000000; assign b = 64'h5F10000000000000;
    #10 assign a = 64'h60CFFFFFFFFFFFFF; assign b = 64'h5F1FFFFFFFFFFFFF;

    #10 $display("\n2**526 * 2**497:");
    #10 assign a = 64'h60D0000000000000; assign b = 64'h5F00000000000000;
    #10 assign a = 64'h60DFFFFFFFFFFFFF; assign b = 64'h5F0FFFFFFFFFFFFF;

    #10 $display("\n2**527 * 2**496:");
    #10 assign a = 64'h60E0000000000000; assign b = 64'h5EF0000000000000;
    #10 assign a = 64'h60EFFFFFFFFFFFFF; assign b = 64'h5EFFFFFFFFFFFFFF;

    #10 $display("\n2**528 * 2**495:");
    #10 assign a = 64'h60F0000000000000; assign b = 64'h5EE0000000000000;
    #10 assign a = 64'h60FFFFFFFFFFFFFF; assign b = 64'h5EEFFFFFFFFFFFFF;

    #10 $display("\n2**529 * 2**494:");
    #10 assign a = 64'h6100000000000000; assign b = 64'h5ED0000000000000;
    #10 assign a = 64'h610FFFFFFFFFFFFF; assign b = 64'h5EDFFFFFFFFFFFFF;

    #10 $display("\n2**530 * 2**493:");
    #10 assign a = 64'h6110000000000000; assign b = 64'h5EC0000000000000;
    #10 assign a = 64'h611FFFFFFFFFFFFF; assign b = 64'h5ECFFFFFFFFFFFFF;

    #10 $display("\n2**531 * 2**492:");
    #10 assign a = 64'h6120000000000000; assign b = 64'h5EB0000000000000;
    #10 assign a = 64'h612FFFFFFFFFFFFF; assign b = 64'h5EBFFFFFFFFFFFFF;

    #10 $display("\n2**532 * 2**491:");
    #10 assign a = 64'h6130000000000000; assign b = 64'h5EA0000000000000;
    #10 assign a = 64'h613FFFFFFFFFFFFF; assign b = 64'h5EAFFFFFFFFFFFFF;

    #10 $display("\n2**533 * 2**490:");
    #10 assign a = 64'h6140000000000000; assign b = 64'h5E90000000000000;
    #10 assign a = 64'h614FFFFFFFFFFFFF; assign b = 64'h5E9FFFFFFFFFFFFF;

    #10 $display("\n2**534 * 2**489:");
    #10 assign a = 64'h6150000000000000; assign b = 64'h5E80000000000000;
    #10 assign a = 64'h615FFFFFFFFFFFFF; assign b = 64'h5E8FFFFFFFFFFFFF;

    #10 $display("\n2**535 * 2**488:");
    #10 assign a = 64'h6160000000000000; assign b = 64'h5E70000000000000;
    #10 assign a = 64'h616FFFFFFFFFFFFF; assign b = 64'h5E7FFFFFFFFFFFFF;

    #10 $display("\n2**536 * 2**487:");
    #10 assign a = 64'h6170000000000000; assign b = 64'h5E60000000000000;
    #10 assign a = 64'h617FFFFFFFFFFFFF; assign b = 64'h5E6FFFFFFFFFFFFF;

    #10 $display("\n2**537 * 2**486:");
    #10 assign a = 64'h6180000000000000; assign b = 64'h5E50000000000000;
    #10 assign a = 64'h618FFFFFFFFFFFFF; assign b = 64'h5E5FFFFFFFFFFFFF;

    #10 $display("\n2**538 * 2**485:");
    #10 assign a = 64'h6190000000000000; assign b = 64'h5E40000000000000;
    #10 assign a = 64'h619FFFFFFFFFFFFF; assign b = 64'h5E4FFFFFFFFFFFFF;

    #10 $display("\n2**539 * 2**484:");
    #10 assign a = 64'h61A0000000000000; assign b = 64'h5E30000000000000;
    #10 assign a = 64'h61AFFFFFFFFFFFFF; assign b = 64'h5E3FFFFFFFFFFFFF;

    #10 $display("\n2**540 * 2**483:");
    #10 assign a = 64'h61B0000000000000; assign b = 64'h5E20000000000000;
    #10 assign a = 64'h61BFFFFFFFFFFFFF; assign b = 64'h5E2FFFFFFFFFFFFF;

    #10 $display("\n2**541 * 2**482:");
    #10 assign a = 64'h61C0000000000000; assign b = 64'h5E10000000000000;
    #10 assign a = 64'h61CFFFFFFFFFFFFF; assign b = 64'h5E1FFFFFFFFFFFFF;

    #10 $display("\n2**542 * 2**481:");
    #10 assign a = 64'h61D0000000000000; assign b = 64'h5E00000000000000;
    #10 assign a = 64'h61DFFFFFFFFFFFFF; assign b = 64'h5E0FFFFFFFFFFFFF;

    #10 $display("\n2**543 * 2**480:");
    #10 assign a = 64'h61E0000000000000; assign b = 64'h5DF0000000000000;
    #10 assign a = 64'h61EFFFFFFFFFFFFF; assign b = 64'h5DFFFFFFFFFFFFFF;

    #10 $display("\n2**544 * 2**479:");
    #10 assign a = 64'h61F0000000000000; assign b = 64'h5DE0000000000000;
    #10 assign a = 64'h61FFFFFFFFFFFFFF; assign b = 64'h5DEFFFFFFFFFFFFF;

    #10 $display("\n2**545 * 2**478:");
    #10 assign a = 64'h6200000000000000; assign b = 64'h5DD0000000000000;
    #10 assign a = 64'h620FFFFFFFFFFFFF; assign b = 64'h5DDFFFFFFFFFFFFF;

    #10 $display("\n2**546 * 2**477:");
    #10 assign a = 64'h6210000000000000; assign b = 64'h5DC0000000000000;
    #10 assign a = 64'h621FFFFFFFFFFFFF; assign b = 64'h5DCFFFFFFFFFFFFF;

    #10 $display("\n2**547 * 2**476:");
    #10 assign a = 64'h6220000000000000; assign b = 64'h5DB0000000000000;
    #10 assign a = 64'h622FFFFFFFFFFFFF; assign b = 64'h5DBFFFFFFFFFFFFF;

    #10 $display("\n2**548 * 2**475:");
    #10 assign a = 64'h6230000000000000; assign b = 64'h5DA0000000000000;
    #10 assign a = 64'h623FFFFFFFFFFFFF; assign b = 64'h5DAFFFFFFFFFFFFF;

    #10 $display("\n2**549 * 2**474:");
    #10 assign a = 64'h6240000000000000; assign b = 64'h5D90000000000000;
    #10 assign a = 64'h624FFFFFFFFFFFFF; assign b = 64'h5D9FFFFFFFFFFFFF;

    #10 $display("\n2**550 * 2**473:");
    #10 assign a = 64'h6250000000000000; assign b = 64'h5D80000000000000;
    #10 assign a = 64'h625FFFFFFFFFFFFF; assign b = 64'h5D8FFFFFFFFFFFFF;

    #10 $display("\n2**551 * 2**472:");
    #10 assign a = 64'h6260000000000000; assign b = 64'h5D70000000000000;
    #10 assign a = 64'h626FFFFFFFFFFFFF; assign b = 64'h5D7FFFFFFFFFFFFF;

    #10 $display("\n2**552 * 2**471:");
    #10 assign a = 64'h6270000000000000; assign b = 64'h5D60000000000000;
    #10 assign a = 64'h627FFFFFFFFFFFFF; assign b = 64'h5D6FFFFFFFFFFFFF;

    #10 $display("\n2**553 * 2**470:");
    #10 assign a = 64'h6280000000000000; assign b = 64'h5D50000000000000;
    #10 assign a = 64'h628FFFFFFFFFFFFF; assign b = 64'h5D5FFFFFFFFFFFFF;

    #10 $display("\n2**554 * 2**469:");
    #10 assign a = 64'h6290000000000000; assign b = 64'h5D40000000000000;
    #10 assign a = 64'h629FFFFFFFFFFFFF; assign b = 64'h5D4FFFFFFFFFFFFF;

    #10 $display("\n2**555 * 2**468:");
    #10 assign a = 64'h62A0000000000000; assign b = 64'h5D30000000000000;
    #10 assign a = 64'h62AFFFFFFFFFFFFF; assign b = 64'h5D3FFFFFFFFFFFFF;

    #10 $display("\n2**556 * 2**467:");
    #10 assign a = 64'h62B0000000000000; assign b = 64'h5D20000000000000;
    #10 assign a = 64'h62BFFFFFFFFFFFFF; assign b = 64'h5D2FFFFFFFFFFFFF;

    #10 $display("\n2**557 * 2**466:");
    #10 assign a = 64'h62C0000000000000; assign b = 64'h5D10000000000000;
    #10 assign a = 64'h62CFFFFFFFFFFFFF; assign b = 64'h5D1FFFFFFFFFFFFF;

    #10 $display("\n2**558 * 2**465:");
    #10 assign a = 64'h62D0000000000000; assign b = 64'h5D00000000000000;
    #10 assign a = 64'h62DFFFFFFFFFFFFF; assign b = 64'h5D0FFFFFFFFFFFFF;

    #10 $display("\n2**559 * 2**464:");
    #10 assign a = 64'h62E0000000000000; assign b = 64'h5CF0000000000000;
    #10 assign a = 64'h62EFFFFFFFFFFFFF; assign b = 64'h5CFFFFFFFFFFFFFF;

    #10 $display("\n2**560 * 2**463:");
    #10 assign a = 64'h62F0000000000000; assign b = 64'h5CE0000000000000;
    #10 assign a = 64'h62FFFFFFFFFFFFFF; assign b = 64'h5CEFFFFFFFFFFFFF;

    #10 $display("\n2**561 * 2**462:");
    #10 assign a = 64'h6300000000000000; assign b = 64'h5CD0000000000000;
    #10 assign a = 64'h630FFFFFFFFFFFFF; assign b = 64'h5CDFFFFFFFFFFFFF;

    #10 $display("\n2**562 * 2**461:");
    #10 assign a = 64'h6310000000000000; assign b = 64'h5CC0000000000000;
    #10 assign a = 64'h631FFFFFFFFFFFFF; assign b = 64'h5CCFFFFFFFFFFFFF;

    #10 $display("\n2**563 * 2**460:");
    #10 assign a = 64'h6320000000000000; assign b = 64'h5CB0000000000000;
    #10 assign a = 64'h632FFFFFFFFFFFFF; assign b = 64'h5CBFFFFFFFFFFFFF;

    #10 $display("\n2**564 * 2**459:");
    #10 assign a = 64'h6330000000000000; assign b = 64'h5CA0000000000000;
    #10 assign a = 64'h633FFFFFFFFFFFFF; assign b = 64'h5CAFFFFFFFFFFFFF;

    #10 $display("\n2**565 * 2**458:");
    #10 assign a = 64'h6340000000000000; assign b = 64'h5C90000000000000;
    #10 assign a = 64'h634FFFFFFFFFFFFF; assign b = 64'h5C9FFFFFFFFFFFFF;

    #10 $display("\n2**566 * 2**457:");
    #10 assign a = 64'h6350000000000000; assign b = 64'h5C80000000000000;
    #10 assign a = 64'h635FFFFFFFFFFFFF; assign b = 64'h5C8FFFFFFFFFFFFF;

    #10 $display("\n2**567 * 2**456:");
    #10 assign a = 64'h6360000000000000; assign b = 64'h5C70000000000000;
    #10 assign a = 64'h636FFFFFFFFFFFFF; assign b = 64'h5C7FFFFFFFFFFFFF;

    #10 $display("\n2**568 * 2**455:");
    #10 assign a = 64'h6370000000000000; assign b = 64'h5C60000000000000;
    #10 assign a = 64'h637FFFFFFFFFFFFF; assign b = 64'h5C6FFFFFFFFFFFFF;

    #10 $display("\n2**569 * 2**454:");
    #10 assign a = 64'h6380000000000000; assign b = 64'h5C50000000000000;
    #10 assign a = 64'h638FFFFFFFFFFFFF; assign b = 64'h5C5FFFFFFFFFFFFF;

    #10 $display("\n2**570 * 2**453:");
    #10 assign a = 64'h6390000000000000; assign b = 64'h5C40000000000000;
    #10 assign a = 64'h639FFFFFFFFFFFFF; assign b = 64'h5C4FFFFFFFFFFFFF;

    #10 $display("\n2**571 * 2**452:");
    #10 assign a = 64'h63A0000000000000; assign b = 64'h5C30000000000000;
    #10 assign a = 64'h63AFFFFFFFFFFFFF; assign b = 64'h5C3FFFFFFFFFFFFF;

    #10 $display("\n2**572 * 2**451:");
    #10 assign a = 64'h63B0000000000000; assign b = 64'h5C20000000000000;
    #10 assign a = 64'h63BFFFFFFFFFFFFF; assign b = 64'h5C2FFFFFFFFFFFFF;

    #10 $display("\n2**573 * 2**450:");
    #10 assign a = 64'h63C0000000000000; assign b = 64'h5C10000000000000;
    #10 assign a = 64'h63CFFFFFFFFFFFFF; assign b = 64'h5C1FFFFFFFFFFFFF;

    #10 $display("\n2**574 * 2**449:");
    #10 assign a = 64'h63D0000000000000; assign b = 64'h5C00000000000000;
    #10 assign a = 64'h63DFFFFFFFFFFFFF; assign b = 64'h5C0FFFFFFFFFFFFF;

    #10 $display("\n2**575 * 2**448:");
    #10 assign a = 64'h63E0000000000000; assign b = 64'h5BF0000000000000;
    #10 assign a = 64'h63EFFFFFFFFFFFFF; assign b = 64'h5BFFFFFFFFFFFFFF;

    #10 $display("\n2**576 * 2**447:");
    #10 assign a = 64'h63F0000000000000; assign b = 64'h5BE0000000000000;
    #10 assign a = 64'h63FFFFFFFFFFFFFF; assign b = 64'h5BEFFFFFFFFFFFFF;

    #10 $display("\n2**577 * 2**446:");
    #10 assign a = 64'h6400000000000000; assign b = 64'h5BD0000000000000;
    #10 assign a = 64'h640FFFFFFFFFFFFF; assign b = 64'h5BDFFFFFFFFFFFFF;

    #10 $display("\n2**578 * 2**445:");
    #10 assign a = 64'h6410000000000000; assign b = 64'h5BC0000000000000;
    #10 assign a = 64'h641FFFFFFFFFFFFF; assign b = 64'h5BCFFFFFFFFFFFFF;

    #10 $display("\n2**579 * 2**444:");
    #10 assign a = 64'h6420000000000000; assign b = 64'h5BB0000000000000;
    #10 assign a = 64'h642FFFFFFFFFFFFF; assign b = 64'h5BBFFFFFFFFFFFFF;

    #10 $display("\n2**580 * 2**443:");
    #10 assign a = 64'h6430000000000000; assign b = 64'h5BA0000000000000;
    #10 assign a = 64'h643FFFFFFFFFFFFF; assign b = 64'h5BAFFFFFFFFFFFFF;

    #10 $display("\n2**581 * 2**442:");
    #10 assign a = 64'h6440000000000000; assign b = 64'h5B90000000000000;
    #10 assign a = 64'h644FFFFFFFFFFFFF; assign b = 64'h5B9FFFFFFFFFFFFF;

    #10 $display("\n2**582 * 2**441:");
    #10 assign a = 64'h6450000000000000; assign b = 64'h5B80000000000000;
    #10 assign a = 64'h645FFFFFFFFFFFFF; assign b = 64'h5B8FFFFFFFFFFFFF;

    #10 $display("\n2**583 * 2**440:");
    #10 assign a = 64'h6460000000000000; assign b = 64'h5B70000000000000;
    #10 assign a = 64'h646FFFFFFFFFFFFF; assign b = 64'h5B7FFFFFFFFFFFFF;

    #10 $display("\n2**584 * 2**439:");
    #10 assign a = 64'h6470000000000000; assign b = 64'h5B60000000000000;
    #10 assign a = 64'h647FFFFFFFFFFFFF; assign b = 64'h5B6FFFFFFFFFFFFF;

    #10 $display("\n2**585 * 2**438:");
    #10 assign a = 64'h6480000000000000; assign b = 64'h5B50000000000000;
    #10 assign a = 64'h648FFFFFFFFFFFFF; assign b = 64'h5B5FFFFFFFFFFFFF;

    #10 $display("\n2**586 * 2**437:");
    #10 assign a = 64'h6490000000000000; assign b = 64'h5B40000000000000;
    #10 assign a = 64'h649FFFFFFFFFFFFF; assign b = 64'h5B4FFFFFFFFFFFFF;

    #10 $display("\n2**587 * 2**436:");
    #10 assign a = 64'h64A0000000000000; assign b = 64'h5B30000000000000;
    #10 assign a = 64'h64AFFFFFFFFFFFFF; assign b = 64'h5B3FFFFFFFFFFFFF;

    #10 $display("\n2**588 * 2**435:");
    #10 assign a = 64'h64B0000000000000; assign b = 64'h5B20000000000000;
    #10 assign a = 64'h64BFFFFFFFFFFFFF; assign b = 64'h5B2FFFFFFFFFFFFF;

    #10 $display("\n2**589 * 2**434:");
    #10 assign a = 64'h64C0000000000000; assign b = 64'h5B10000000000000;
    #10 assign a = 64'h64CFFFFFFFFFFFFF; assign b = 64'h5B1FFFFFFFFFFFFF;

    #10 $display("\n2**590 * 2**433:");
    #10 assign a = 64'h64D0000000000000; assign b = 64'h5B00000000000000;
    #10 assign a = 64'h64DFFFFFFFFFFFFF; assign b = 64'h5B0FFFFFFFFFFFFF;

    #10 $display("\n2**591 * 2**432:");
    #10 assign a = 64'h64E0000000000000; assign b = 64'h5AF0000000000000;
    #10 assign a = 64'h64EFFFFFFFFFFFFF; assign b = 64'h5AFFFFFFFFFFFFFF;

    #10 $display("\n2**592 * 2**431:");
    #10 assign a = 64'h64F0000000000000; assign b = 64'h5AE0000000000000;
    #10 assign a = 64'h64FFFFFFFFFFFFFF; assign b = 64'h5AEFFFFFFFFFFFFF;

    #10 $display("\n2**593 * 2**430:");
    #10 assign a = 64'h6500000000000000; assign b = 64'h5AD0000000000000;
    #10 assign a = 64'h650FFFFFFFFFFFFF; assign b = 64'h5ADFFFFFFFFFFFFF;

    #10 $display("\n2**594 * 2**429:");
    #10 assign a = 64'h6510000000000000; assign b = 64'h5AC0000000000000;
    #10 assign a = 64'h651FFFFFFFFFFFFF; assign b = 64'h5ACFFFFFFFFFFFFF;

    #10 $display("\n2**595 * 2**428:");
    #10 assign a = 64'h6520000000000000; assign b = 64'h5AB0000000000000;
    #10 assign a = 64'h652FFFFFFFFFFFFF; assign b = 64'h5ABFFFFFFFFFFFFF;

    #10 $display("\n2**596 * 2**427:");
    #10 assign a = 64'h6530000000000000; assign b = 64'h5AA0000000000000;
    #10 assign a = 64'h653FFFFFFFFFFFFF; assign b = 64'h5AAFFFFFFFFFFFFF;

    #10 $display("\n2**597 * 2**426:");
    #10 assign a = 64'h6540000000000000; assign b = 64'h5A90000000000000;
    #10 assign a = 64'h654FFFFFFFFFFFFF; assign b = 64'h5A9FFFFFFFFFFFFF;

    #10 $display("\n2**598 * 2**425:");
    #10 assign a = 64'h6550000000000000; assign b = 64'h5A80000000000000;
    #10 assign a = 64'h655FFFFFFFFFFFFF; assign b = 64'h5A8FFFFFFFFFFFFF;

    #10 $display("\n2**599 * 2**424:");
    #10 assign a = 64'h6560000000000000; assign b = 64'h5A70000000000000;
    #10 assign a = 64'h656FFFFFFFFFFFFF; assign b = 64'h5A7FFFFFFFFFFFFF;

    #10 $display("\n2**600 * 2**423:");
    #10 assign a = 64'h6570000000000000; assign b = 64'h5A60000000000000;
    #10 assign a = 64'h657FFFFFFFFFFFFF; assign b = 64'h5A6FFFFFFFFFFFFF;

    #10 $display("\n2**601 * 2**422:");
    #10 assign a = 64'h6580000000000000; assign b = 64'h5A50000000000000;
    #10 assign a = 64'h658FFFFFFFFFFFFF; assign b = 64'h5A5FFFFFFFFFFFFF;

    #10 $display("\n2**602 * 2**421:");
    #10 assign a = 64'h6590000000000000; assign b = 64'h5A40000000000000;
    #10 assign a = 64'h659FFFFFFFFFFFFF; assign b = 64'h5A4FFFFFFFFFFFFF;

    #10 $display("\n2**603 * 2**420:");
    #10 assign a = 64'h65A0000000000000; assign b = 64'h5A30000000000000;
    #10 assign a = 64'h65AFFFFFFFFFFFFF; assign b = 64'h5A3FFFFFFFFFFFFF;

    #10 $display("\n2**604 * 2**419:");
    #10 assign a = 64'h65B0000000000000; assign b = 64'h5A20000000000000;
    #10 assign a = 64'h65BFFFFFFFFFFFFF; assign b = 64'h5A2FFFFFFFFFFFFF;

    #10 $display("\n2**605 * 2**418:");
    #10 assign a = 64'h65C0000000000000; assign b = 64'h5A10000000000000;
    #10 assign a = 64'h65CFFFFFFFFFFFFF; assign b = 64'h5A1FFFFFFFFFFFFF;

    #10 $display("\n2**606 * 2**417:");
    #10 assign a = 64'h65D0000000000000; assign b = 64'h5A00000000000000;
    #10 assign a = 64'h65DFFFFFFFFFFFFF; assign b = 64'h5A0FFFFFFFFFFFFF;

    #10 $display("\n2**607 * 2**416:");
    #10 assign a = 64'h65E0000000000000; assign b = 64'h59F0000000000000;
    #10 assign a = 64'h65EFFFFFFFFFFFFF; assign b = 64'h59FFFFFFFFFFFFFF;

    #10 $display("\n2**608 * 2**415:");
    #10 assign a = 64'h65F0000000000000; assign b = 64'h59E0000000000000;
    #10 assign a = 64'h65FFFFFFFFFFFFFF; assign b = 64'h59EFFFFFFFFFFFFF;

    #10 $display("\n2**609 * 2**414:");
    #10 assign a = 64'h6600000000000000; assign b = 64'h59D0000000000000;
    #10 assign a = 64'h660FFFFFFFFFFFFF; assign b = 64'h59DFFFFFFFFFFFFF;

    #10 $display("\n2**610 * 2**413:");
    #10 assign a = 64'h6610000000000000; assign b = 64'h59C0000000000000;
    #10 assign a = 64'h661FFFFFFFFFFFFF; assign b = 64'h59CFFFFFFFFFFFFF;

    #10 $display("\n2**611 * 2**412:");
    #10 assign a = 64'h6620000000000000; assign b = 64'h59B0000000000000;
    #10 assign a = 64'h662FFFFFFFFFFFFF; assign b = 64'h59BFFFFFFFFFFFFF;

    #10 $display("\n2**612 * 2**411:");
    #10 assign a = 64'h6630000000000000; assign b = 64'h59A0000000000000;
    #10 assign a = 64'h663FFFFFFFFFFFFF; assign b = 64'h59AFFFFFFFFFFFFF;

    #10 $display("\n2**613 * 2**410:");
    #10 assign a = 64'h6640000000000000; assign b = 64'h5990000000000000;
    #10 assign a = 64'h664FFFFFFFFFFFFF; assign b = 64'h599FFFFFFFFFFFFF;

    #10 $display("\n2**614 * 2**409:");
    #10 assign a = 64'h6650000000000000; assign b = 64'h5980000000000000;
    #10 assign a = 64'h665FFFFFFFFFFFFF; assign b = 64'h598FFFFFFFFFFFFF;

    #10 $display("\n2**615 * 2**408:");
    #10 assign a = 64'h6660000000000000; assign b = 64'h5970000000000000;
    #10 assign a = 64'h666FFFFFFFFFFFFF; assign b = 64'h597FFFFFFFFFFFFF;

    #10 $display("\n2**616 * 2**407:");
    #10 assign a = 64'h6670000000000000; assign b = 64'h5960000000000000;
    #10 assign a = 64'h667FFFFFFFFFFFFF; assign b = 64'h596FFFFFFFFFFFFF;

    #10 $display("\n2**617 * 2**406:");
    #10 assign a = 64'h6680000000000000; assign b = 64'h5950000000000000;
    #10 assign a = 64'h668FFFFFFFFFFFFF; assign b = 64'h595FFFFFFFFFFFFF;

    #10 $display("\n2**618 * 2**405:");
    #10 assign a = 64'h6690000000000000; assign b = 64'h5940000000000000;
    #10 assign a = 64'h669FFFFFFFFFFFFF; assign b = 64'h594FFFFFFFFFFFFF;

    #10 $display("\n2**619 * 2**404:");
    #10 assign a = 64'h66A0000000000000; assign b = 64'h5930000000000000;
    #10 assign a = 64'h66AFFFFFFFFFFFFF; assign b = 64'h593FFFFFFFFFFFFF;

    #10 $display("\n2**620 * 2**403:");
    #10 assign a = 64'h66B0000000000000; assign b = 64'h5920000000000000;
    #10 assign a = 64'h66BFFFFFFFFFFFFF; assign b = 64'h592FFFFFFFFFFFFF;

    #10 $display("\n2**621 * 2**402:");
    #10 assign a = 64'h66C0000000000000; assign b = 64'h5910000000000000;
    #10 assign a = 64'h66CFFFFFFFFFFFFF; assign b = 64'h591FFFFFFFFFFFFF;

    #10 $display("\n2**622 * 2**401:");
    #10 assign a = 64'h66D0000000000000; assign b = 64'h5900000000000000;
    #10 assign a = 64'h66DFFFFFFFFFFFFF; assign b = 64'h590FFFFFFFFFFFFF;

    #10 $display("\n2**623 * 2**400:");
    #10 assign a = 64'h66E0000000000000; assign b = 64'h58F0000000000000;
    #10 assign a = 64'h66EFFFFFFFFFFFFF; assign b = 64'h58FFFFFFFFFFFFFF;

    #10 $display("\n2**624 * 2**399:");
    #10 assign a = 64'h66F0000000000000; assign b = 64'h58E0000000000000;
    #10 assign a = 64'h66FFFFFFFFFFFFFF; assign b = 64'h58EFFFFFFFFFFFFF;

    #10 $display("\n2**625 * 2**398:");
    #10 assign a = 64'h6700000000000000; assign b = 64'h58D0000000000000;
    #10 assign a = 64'h670FFFFFFFFFFFFF; assign b = 64'h58DFFFFFFFFFFFFF;

    #10 $display("\n2**626 * 2**397:");
    #10 assign a = 64'h6710000000000000; assign b = 64'h58C0000000000000;
    #10 assign a = 64'h671FFFFFFFFFFFFF; assign b = 64'h58CFFFFFFFFFFFFF;

    #10 $display("\n2**627 * 2**396:");
    #10 assign a = 64'h6720000000000000; assign b = 64'h58B0000000000000;
    #10 assign a = 64'h672FFFFFFFFFFFFF; assign b = 64'h58BFFFFFFFFFFFFF;

    #10 $display("\n2**628 * 2**395:");
    #10 assign a = 64'h6730000000000000; assign b = 64'h58A0000000000000;
    #10 assign a = 64'h673FFFFFFFFFFFFF; assign b = 64'h58AFFFFFFFFFFFFF;

    #10 $display("\n2**629 * 2**394:");
    #10 assign a = 64'h6740000000000000; assign b = 64'h5890000000000000;
    #10 assign a = 64'h674FFFFFFFFFFFFF; assign b = 64'h589FFFFFFFFFFFFF;

    #10 $display("\n2**630 * 2**393:");
    #10 assign a = 64'h6750000000000000; assign b = 64'h5880000000000000;
    #10 assign a = 64'h675FFFFFFFFFFFFF; assign b = 64'h588FFFFFFFFFFFFF;

    #10 $display("\n2**631 * 2**392:");
    #10 assign a = 64'h6760000000000000; assign b = 64'h5870000000000000;
    #10 assign a = 64'h676FFFFFFFFFFFFF; assign b = 64'h587FFFFFFFFFFFFF;

    #10 $display("\n2**632 * 2**391:");
    #10 assign a = 64'h6770000000000000; assign b = 64'h5860000000000000;
    #10 assign a = 64'h677FFFFFFFFFFFFF; assign b = 64'h586FFFFFFFFFFFFF;

    #10 $display("\n2**633 * 2**390:");
    #10 assign a = 64'h6780000000000000; assign b = 64'h5850000000000000;
    #10 assign a = 64'h678FFFFFFFFFFFFF; assign b = 64'h585FFFFFFFFFFFFF;

    #10 $display("\n2**634 * 2**389:");
    #10 assign a = 64'h6790000000000000; assign b = 64'h5840000000000000;
    #10 assign a = 64'h679FFFFFFFFFFFFF; assign b = 64'h584FFFFFFFFFFFFF;

    #10 $display("\n2**635 * 2**388:");
    #10 assign a = 64'h67A0000000000000; assign b = 64'h5830000000000000;
    #10 assign a = 64'h67AFFFFFFFFFFFFF; assign b = 64'h583FFFFFFFFFFFFF;

    #10 $display("\n2**636 * 2**387:");
    #10 assign a = 64'h67B0000000000000; assign b = 64'h5820000000000000;
    #10 assign a = 64'h67BFFFFFFFFFFFFF; assign b = 64'h582FFFFFFFFFFFFF;

    #10 $display("\n2**637 * 2**386:");
    #10 assign a = 64'h67C0000000000000; assign b = 64'h5810000000000000;
    #10 assign a = 64'h67CFFFFFFFFFFFFF; assign b = 64'h581FFFFFFFFFFFFF;

    #10 $display("\n2**638 * 2**385:");
    #10 assign a = 64'h67D0000000000000; assign b = 64'h5800000000000000;
    #10 assign a = 64'h67DFFFFFFFFFFFFF; assign b = 64'h580FFFFFFFFFFFFF;

    #10 $display("\n2**639 * 2**384:");
    #10 assign a = 64'h67E0000000000000; assign b = 64'h57F0000000000000;
    #10 assign a = 64'h67EFFFFFFFFFFFFF; assign b = 64'h57FFFFFFFFFFFFFF;

    #10 $display("\n2**640 * 2**383:");
    #10 assign a = 64'h67F0000000000000; assign b = 64'h57E0000000000000;
    #10 assign a = 64'h67FFFFFFFFFFFFFF; assign b = 64'h57EFFFFFFFFFFFFF;

    #10 $display("\n2**641 * 2**382:");
    #10 assign a = 64'h6800000000000000; assign b = 64'h57D0000000000000;
    #10 assign a = 64'h680FFFFFFFFFFFFF; assign b = 64'h57DFFFFFFFFFFFFF;

    #10 $display("\n2**642 * 2**381:");
    #10 assign a = 64'h6810000000000000; assign b = 64'h57C0000000000000;
    #10 assign a = 64'h681FFFFFFFFFFFFF; assign b = 64'h57CFFFFFFFFFFFFF;

    #10 $display("\n2**643 * 2**380:");
    #10 assign a = 64'h6820000000000000; assign b = 64'h57B0000000000000;
    #10 assign a = 64'h682FFFFFFFFFFFFF; assign b = 64'h57BFFFFFFFFFFFFF;

    #10 $display("\n2**644 * 2**379:");
    #10 assign a = 64'h6830000000000000; assign b = 64'h57A0000000000000;
    #10 assign a = 64'h683FFFFFFFFFFFFF; assign b = 64'h57AFFFFFFFFFFFFF;

    #10 $display("\n2**645 * 2**378:");
    #10 assign a = 64'h6840000000000000; assign b = 64'h5790000000000000;
    #10 assign a = 64'h684FFFFFFFFFFFFF; assign b = 64'h579FFFFFFFFFFFFF;

    #10 $display("\n2**646 * 2**377:");
    #10 assign a = 64'h6850000000000000; assign b = 64'h5780000000000000;
    #10 assign a = 64'h685FFFFFFFFFFFFF; assign b = 64'h578FFFFFFFFFFFFF;

    #10 $display("\n2**647 * 2**376:");
    #10 assign a = 64'h6860000000000000; assign b = 64'h5770000000000000;
    #10 assign a = 64'h686FFFFFFFFFFFFF; assign b = 64'h577FFFFFFFFFFFFF;

    #10 $display("\n2**648 * 2**375:");
    #10 assign a = 64'h6870000000000000; assign b = 64'h5760000000000000;
    #10 assign a = 64'h687FFFFFFFFFFFFF; assign b = 64'h576FFFFFFFFFFFFF;

    #10 $display("\n2**649 * 2**374:");
    #10 assign a = 64'h6880000000000000; assign b = 64'h5750000000000000;
    #10 assign a = 64'h688FFFFFFFFFFFFF; assign b = 64'h575FFFFFFFFFFFFF;

    #10 $display("\n2**650 * 2**373:");
    #10 assign a = 64'h6890000000000000; assign b = 64'h5740000000000000;
    #10 assign a = 64'h689FFFFFFFFFFFFF; assign b = 64'h574FFFFFFFFFFFFF;

    #10 $display("\n2**651 * 2**372:");
    #10 assign a = 64'h68A0000000000000; assign b = 64'h5730000000000000;
    #10 assign a = 64'h68AFFFFFFFFFFFFF; assign b = 64'h573FFFFFFFFFFFFF;

    #10 $display("\n2**652 * 2**371:");
    #10 assign a = 64'h68B0000000000000; assign b = 64'h5720000000000000;
    #10 assign a = 64'h68BFFFFFFFFFFFFF; assign b = 64'h572FFFFFFFFFFFFF;

    #10 $display("\n2**653 * 2**370:");
    #10 assign a = 64'h68C0000000000000; assign b = 64'h5710000000000000;
    #10 assign a = 64'h68CFFFFFFFFFFFFF; assign b = 64'h571FFFFFFFFFFFFF;

    #10 $display("\n2**654 * 2**369:");
    #10 assign a = 64'h68D0000000000000; assign b = 64'h5700000000000000;
    #10 assign a = 64'h68DFFFFFFFFFFFFF; assign b = 64'h570FFFFFFFFFFFFF;

    #10 $display("\n2**655 * 2**368:");
    #10 assign a = 64'h68E0000000000000; assign b = 64'h56F0000000000000;
    #10 assign a = 64'h68EFFFFFFFFFFFFF; assign b = 64'h56FFFFFFFFFFFFFF;

    #10 $display("\n2**656 * 2**367:");
    #10 assign a = 64'h68F0000000000000; assign b = 64'h56E0000000000000;
    #10 assign a = 64'h68FFFFFFFFFFFFFF; assign b = 64'h56EFFFFFFFFFFFFF;

    #10 $display("\n2**657 * 2**366:");
    #10 assign a = 64'h6900000000000000; assign b = 64'h56D0000000000000;
    #10 assign a = 64'h690FFFFFFFFFFFFF; assign b = 64'h56DFFFFFFFFFFFFF;

    #10 $display("\n2**658 * 2**365:");
    #10 assign a = 64'h6910000000000000; assign b = 64'h56C0000000000000;
    #10 assign a = 64'h691FFFFFFFFFFFFF; assign b = 64'h56CFFFFFFFFFFFFF;

    #10 $display("\n2**659 * 2**364:");
    #10 assign a = 64'h6920000000000000; assign b = 64'h56B0000000000000;
    #10 assign a = 64'h692FFFFFFFFFFFFF; assign b = 64'h56BFFFFFFFFFFFFF;

    #10 $display("\n2**660 * 2**363:");
    #10 assign a = 64'h6930000000000000; assign b = 64'h56A0000000000000;
    #10 assign a = 64'h693FFFFFFFFFFFFF; assign b = 64'h56AFFFFFFFFFFFFF;

    #10 $display("\n2**661 * 2**362:");
    #10 assign a = 64'h6940000000000000; assign b = 64'h5690000000000000;
    #10 assign a = 64'h694FFFFFFFFFFFFF; assign b = 64'h569FFFFFFFFFFFFF;

    #10 $display("\n2**662 * 2**361:");
    #10 assign a = 64'h6950000000000000; assign b = 64'h5680000000000000;
    #10 assign a = 64'h695FFFFFFFFFFFFF; assign b = 64'h568FFFFFFFFFFFFF;

    #10 $display("\n2**663 * 2**360:");
    #10 assign a = 64'h6960000000000000; assign b = 64'h5670000000000000;
    #10 assign a = 64'h696FFFFFFFFFFFFF; assign b = 64'h567FFFFFFFFFFFFF;

    #10 $display("\n2**664 * 2**359:");
    #10 assign a = 64'h6970000000000000; assign b = 64'h5660000000000000;
    #10 assign a = 64'h697FFFFFFFFFFFFF; assign b = 64'h566FFFFFFFFFFFFF;

    #10 $display("\n2**665 * 2**358:");
    #10 assign a = 64'h6980000000000000; assign b = 64'h5650000000000000;
    #10 assign a = 64'h698FFFFFFFFFFFFF; assign b = 64'h565FFFFFFFFFFFFF;

    #10 $display("\n2**666 * 2**357:");
    #10 assign a = 64'h6990000000000000; assign b = 64'h5640000000000000;
    #10 assign a = 64'h699FFFFFFFFFFFFF; assign b = 64'h564FFFFFFFFFFFFF;

    #10 $display("\n2**667 * 2**356:");
    #10 assign a = 64'h69A0000000000000; assign b = 64'h5630000000000000;
    #10 assign a = 64'h69AFFFFFFFFFFFFF; assign b = 64'h563FFFFFFFFFFFFF;

    #10 $display("\n2**668 * 2**355:");
    #10 assign a = 64'h69B0000000000000; assign b = 64'h5620000000000000;
    #10 assign a = 64'h69BFFFFFFFFFFFFF; assign b = 64'h562FFFFFFFFFFFFF;

    #10 $display("\n2**669 * 2**354:");
    #10 assign a = 64'h69C0000000000000; assign b = 64'h5610000000000000;
    #10 assign a = 64'h69CFFFFFFFFFFFFF; assign b = 64'h561FFFFFFFFFFFFF;

    #10 $display("\n2**670 * 2**353:");
    #10 assign a = 64'h69D0000000000000; assign b = 64'h5600000000000000;
    #10 assign a = 64'h69DFFFFFFFFFFFFF; assign b = 64'h560FFFFFFFFFFFFF;

    #10 $display("\n2**671 * 2**352:");
    #10 assign a = 64'h69E0000000000000; assign b = 64'h55F0000000000000;
    #10 assign a = 64'h69EFFFFFFFFFFFFF; assign b = 64'h55FFFFFFFFFFFFFF;

    #10 $display("\n2**672 * 2**351:");
    #10 assign a = 64'h69F0000000000000; assign b = 64'h55E0000000000000;
    #10 assign a = 64'h69FFFFFFFFFFFFFF; assign b = 64'h55EFFFFFFFFFFFFF;

    #10 $display("\n2**673 * 2**350:");
    #10 assign a = 64'h6A00000000000000; assign b = 64'h55D0000000000000;
    #10 assign a = 64'h6A0FFFFFFFFFFFFF; assign b = 64'h55DFFFFFFFFFFFFF;

    #10 $display("\n2**674 * 2**349:");
    #10 assign a = 64'h6A10000000000000; assign b = 64'h55C0000000000000;
    #10 assign a = 64'h6A1FFFFFFFFFFFFF; assign b = 64'h55CFFFFFFFFFFFFF;

    #10 $display("\n2**675 * 2**348:");
    #10 assign a = 64'h6A20000000000000; assign b = 64'h55B0000000000000;
    #10 assign a = 64'h6A2FFFFFFFFFFFFF; assign b = 64'h55BFFFFFFFFFFFFF;

    #10 $display("\n2**676 * 2**347:");
    #10 assign a = 64'h6A30000000000000; assign b = 64'h55A0000000000000;
    #10 assign a = 64'h6A3FFFFFFFFFFFFF; assign b = 64'h55AFFFFFFFFFFFFF;

    #10 $display("\n2**677 * 2**346:");
    #10 assign a = 64'h6A40000000000000; assign b = 64'h5590000000000000;
    #10 assign a = 64'h6A4FFFFFFFFFFFFF; assign b = 64'h559FFFFFFFFFFFFF;

    #10 $display("\n2**678 * 2**345:");
    #10 assign a = 64'h6A50000000000000; assign b = 64'h5580000000000000;
    #10 assign a = 64'h6A5FFFFFFFFFFFFF; assign b = 64'h558FFFFFFFFFFFFF;

    #10 $display("\n2**679 * 2**344:");
    #10 assign a = 64'h6A60000000000000; assign b = 64'h5570000000000000;
    #10 assign a = 64'h6A6FFFFFFFFFFFFF; assign b = 64'h557FFFFFFFFFFFFF;

    #10 $display("\n2**680 * 2**343:");
    #10 assign a = 64'h6A70000000000000; assign b = 64'h5560000000000000;
    #10 assign a = 64'h6A7FFFFFFFFFFFFF; assign b = 64'h556FFFFFFFFFFFFF;

    #10 $display("\n2**681 * 2**342:");
    #10 assign a = 64'h6A80000000000000; assign b = 64'h5550000000000000;
    #10 assign a = 64'h6A8FFFFFFFFFFFFF; assign b = 64'h555FFFFFFFFFFFFF;

    #10 $display("\n2**682 * 2**341:");
    #10 assign a = 64'h6A90000000000000; assign b = 64'h5540000000000000;
    #10 assign a = 64'h6A9FFFFFFFFFFFFF; assign b = 64'h554FFFFFFFFFFFFF;

    #10 $display("\n2**683 * 2**340:");
    #10 assign a = 64'h6AA0000000000000; assign b = 64'h5530000000000000;
    #10 assign a = 64'h6AAFFFFFFFFFFFFF; assign b = 64'h553FFFFFFFFFFFFF;

    #10 $display("\n2**684 * 2**339:");
    #10 assign a = 64'h6AB0000000000000; assign b = 64'h5520000000000000;
    #10 assign a = 64'h6ABFFFFFFFFFFFFF; assign b = 64'h552FFFFFFFFFFFFF;

    #10 $display("\n2**685 * 2**338:");
    #10 assign a = 64'h6AC0000000000000; assign b = 64'h5510000000000000;
    #10 assign a = 64'h6ACFFFFFFFFFFFFF; assign b = 64'h551FFFFFFFFFFFFF;

    #10 $display("\n2**686 * 2**337:");
    #10 assign a = 64'h6AD0000000000000; assign b = 64'h5500000000000000;
    #10 assign a = 64'h6ADFFFFFFFFFFFFF; assign b = 64'h550FFFFFFFFFFFFF;

    #10 $display("\n2**687 * 2**336:");
    #10 assign a = 64'h6AE0000000000000; assign b = 64'h54F0000000000000;
    #10 assign a = 64'h6AEFFFFFFFFFFFFF; assign b = 64'h54FFFFFFFFFFFFFF;

    #10 $display("\n2**688 * 2**335:");
    #10 assign a = 64'h6AF0000000000000; assign b = 64'h54E0000000000000;
    #10 assign a = 64'h6AFFFFFFFFFFFFFF; assign b = 64'h54EFFFFFFFFFFFFF;

    #10 $display("\n2**689 * 2**334:");
    #10 assign a = 64'h6B00000000000000; assign b = 64'h54D0000000000000;
    #10 assign a = 64'h6B0FFFFFFFFFFFFF; assign b = 64'h54DFFFFFFFFFFFFF;

    #10 $display("\n2**690 * 2**333:");
    #10 assign a = 64'h6B10000000000000; assign b = 64'h54C0000000000000;
    #10 assign a = 64'h6B1FFFFFFFFFFFFF; assign b = 64'h54CFFFFFFFFFFFFF;

    #10 $display("\n2**691 * 2**332:");
    #10 assign a = 64'h6B20000000000000; assign b = 64'h54B0000000000000;
    #10 assign a = 64'h6B2FFFFFFFFFFFFF; assign b = 64'h54BFFFFFFFFFFFFF;

    #10 $display("\n2**692 * 2**331:");
    #10 assign a = 64'h6B30000000000000; assign b = 64'h54A0000000000000;
    #10 assign a = 64'h6B3FFFFFFFFFFFFF; assign b = 64'h54AFFFFFFFFFFFFF;

    #10 $display("\n2**693 * 2**330:");
    #10 assign a = 64'h6B40000000000000; assign b = 64'h5490000000000000;
    #10 assign a = 64'h6B4FFFFFFFFFFFFF; assign b = 64'h549FFFFFFFFFFFFF;

    #10 $display("\n2**694 * 2**329:");
    #10 assign a = 64'h6B50000000000000; assign b = 64'h5480000000000000;
    #10 assign a = 64'h6B5FFFFFFFFFFFFF; assign b = 64'h548FFFFFFFFFFFFF;

    #10 $display("\n2**695 * 2**328:");
    #10 assign a = 64'h6B60000000000000; assign b = 64'h5470000000000000;
    #10 assign a = 64'h6B6FFFFFFFFFFFFF; assign b = 64'h547FFFFFFFFFFFFF;

    #10 $display("\n2**696 * 2**327:");
    #10 assign a = 64'h6B70000000000000; assign b = 64'h5460000000000000;
    #10 assign a = 64'h6B7FFFFFFFFFFFFF; assign b = 64'h546FFFFFFFFFFFFF;

    #10 $display("\n2**697 * 2**326:");
    #10 assign a = 64'h6B80000000000000; assign b = 64'h5450000000000000;
    #10 assign a = 64'h6B8FFFFFFFFFFFFF; assign b = 64'h545FFFFFFFFFFFFF;

    #10 $display("\n2**698 * 2**325:");
    #10 assign a = 64'h6B90000000000000; assign b = 64'h5440000000000000;
    #10 assign a = 64'h6B9FFFFFFFFFFFFF; assign b = 64'h544FFFFFFFFFFFFF;

    #10 $display("\n2**699 * 2**324:");
    #10 assign a = 64'h6BA0000000000000; assign b = 64'h5430000000000000;
    #10 assign a = 64'h6BAFFFFFFFFFFFFF; assign b = 64'h543FFFFFFFFFFFFF;

    #10 $display("\n2**700 * 2**323:");
    #10 assign a = 64'h6BB0000000000000; assign b = 64'h5420000000000000;
    #10 assign a = 64'h6BBFFFFFFFFFFFFF; assign b = 64'h542FFFFFFFFFFFFF;

    #10 $display("\n2**701 * 2**322:");
    #10 assign a = 64'h6BC0000000000000; assign b = 64'h5410000000000000;
    #10 assign a = 64'h6BCFFFFFFFFFFFFF; assign b = 64'h541FFFFFFFFFFFFF;

    #10 $display("\n2**702 * 2**321:");
    #10 assign a = 64'h6BD0000000000000; assign b = 64'h5400000000000000;
    #10 assign a = 64'h6BDFFFFFFFFFFFFF; assign b = 64'h540FFFFFFFFFFFFF;

    #10 $display("\n2**703 * 2**320:");
    #10 assign a = 64'h6BE0000000000000; assign b = 64'h53F0000000000000;
    #10 assign a = 64'h6BEFFFFFFFFFFFFF; assign b = 64'h53FFFFFFFFFFFFFF;

    #10 $display("\n2**704 * 2**319:");
    #10 assign a = 64'h6BF0000000000000; assign b = 64'h53E0000000000000;
    #10 assign a = 64'h6BFFFFFFFFFFFFFF; assign b = 64'h53EFFFFFFFFFFFFF;

    #10 $display("\n2**705 * 2**318:");
    #10 assign a = 64'h6C00000000000000; assign b = 64'h53D0000000000000;
    #10 assign a = 64'h6C0FFFFFFFFFFFFF; assign b = 64'h53DFFFFFFFFFFFFF;

    #10 $display("\n2**706 * 2**317:");
    #10 assign a = 64'h6C10000000000000; assign b = 64'h53C0000000000000;
    #10 assign a = 64'h6C1FFFFFFFFFFFFF; assign b = 64'h53CFFFFFFFFFFFFF;

    #10 $display("\n2**707 * 2**316:");
    #10 assign a = 64'h6C20000000000000; assign b = 64'h53B0000000000000;
    #10 assign a = 64'h6C2FFFFFFFFFFFFF; assign b = 64'h53BFFFFFFFFFFFFF;

    #10 $display("\n2**708 * 2**315:");
    #10 assign a = 64'h6C30000000000000; assign b = 64'h53A0000000000000;
    #10 assign a = 64'h6C3FFFFFFFFFFFFF; assign b = 64'h53AFFFFFFFFFFFFF;

    #10 $display("\n2**709 * 2**314:");
    #10 assign a = 64'h6C40000000000000; assign b = 64'h5390000000000000;
    #10 assign a = 64'h6C4FFFFFFFFFFFFF; assign b = 64'h539FFFFFFFFFFFFF;

    #10 $display("\n2**710 * 2**313:");
    #10 assign a = 64'h6C50000000000000; assign b = 64'h5380000000000000;
    #10 assign a = 64'h6C5FFFFFFFFFFFFF; assign b = 64'h538FFFFFFFFFFFFF;

    #10 $display("\n2**711 * 2**312:");
    #10 assign a = 64'h6C60000000000000; assign b = 64'h5370000000000000;
    #10 assign a = 64'h6C6FFFFFFFFFFFFF; assign b = 64'h537FFFFFFFFFFFFF;

    #10 $display("\n2**712 * 2**311:");
    #10 assign a = 64'h6C70000000000000; assign b = 64'h5360000000000000;
    #10 assign a = 64'h6C7FFFFFFFFFFFFF; assign b = 64'h536FFFFFFFFFFFFF;

    #10 $display("\n2**713 * 2**310:");
    #10 assign a = 64'h6C80000000000000; assign b = 64'h5350000000000000;
    #10 assign a = 64'h6C8FFFFFFFFFFFFF; assign b = 64'h535FFFFFFFFFFFFF;

    #10 $display("\n2**714 * 2**309:");
    #10 assign a = 64'h6C90000000000000; assign b = 64'h5340000000000000;
    #10 assign a = 64'h6C9FFFFFFFFFFFFF; assign b = 64'h534FFFFFFFFFFFFF;

    #10 $display("\n2**715 * 2**308:");
    #10 assign a = 64'h6CA0000000000000; assign b = 64'h5330000000000000;
    #10 assign a = 64'h6CAFFFFFFFFFFFFF; assign b = 64'h533FFFFFFFFFFFFF;

    #10 $display("\n2**716 * 2**307:");
    #10 assign a = 64'h6CB0000000000000; assign b = 64'h5320000000000000;
    #10 assign a = 64'h6CBFFFFFFFFFFFFF; assign b = 64'h532FFFFFFFFFFFFF;

    #10 $display("\n2**717 * 2**306:");
    #10 assign a = 64'h6CC0000000000000; assign b = 64'h5310000000000000;
    #10 assign a = 64'h6CCFFFFFFFFFFFFF; assign b = 64'h531FFFFFFFFFFFFF;

    #10 $display("\n2**718 * 2**305:");
    #10 assign a = 64'h6CD0000000000000; assign b = 64'h5300000000000000;
    #10 assign a = 64'h6CDFFFFFFFFFFFFF; assign b = 64'h530FFFFFFFFFFFFF;

    #10 $display("\n2**719 * 2**304:");
    #10 assign a = 64'h6CE0000000000000; assign b = 64'h52F0000000000000;
    #10 assign a = 64'h6CEFFFFFFFFFFFFF; assign b = 64'h52FFFFFFFFFFFFFF;

    #10 $display("\n2**720 * 2**303:");
    #10 assign a = 64'h6CF0000000000000; assign b = 64'h52E0000000000000;
    #10 assign a = 64'h6CFFFFFFFFFFFFFF; assign b = 64'h52EFFFFFFFFFFFFF;

    #10 $display("\n2**721 * 2**302:");
    #10 assign a = 64'h6D00000000000000; assign b = 64'h52D0000000000000;
    #10 assign a = 64'h6D0FFFFFFFFFFFFF; assign b = 64'h52DFFFFFFFFFFFFF;

    #10 $display("\n2**722 * 2**301:");
    #10 assign a = 64'h6D10000000000000; assign b = 64'h52C0000000000000;
    #10 assign a = 64'h6D1FFFFFFFFFFFFF; assign b = 64'h52CFFFFFFFFFFFFF;

    #10 $display("\n2**723 * 2**300:");
    #10 assign a = 64'h6D20000000000000; assign b = 64'h52B0000000000000;
    #10 assign a = 64'h6D2FFFFFFFFFFFFF; assign b = 64'h52BFFFFFFFFFFFFF;

    #10 $display("\n2**724 * 2**299:");
    #10 assign a = 64'h6D30000000000000; assign b = 64'h52A0000000000000;
    #10 assign a = 64'h6D3FFFFFFFFFFFFF; assign b = 64'h52AFFFFFFFFFFFFF;

    #10 $display("\n2**725 * 2**298:");
    #10 assign a = 64'h6D40000000000000; assign b = 64'h5290000000000000;
    #10 assign a = 64'h6D4FFFFFFFFFFFFF; assign b = 64'h529FFFFFFFFFFFFF;

    #10 $display("\n2**726 * 2**297:");
    #10 assign a = 64'h6D50000000000000; assign b = 64'h5280000000000000;
    #10 assign a = 64'h6D5FFFFFFFFFFFFF; assign b = 64'h528FFFFFFFFFFFFF;

    #10 $display("\n2**727 * 2**296:");
    #10 assign a = 64'h6D60000000000000; assign b = 64'h5270000000000000;
    #10 assign a = 64'h6D6FFFFFFFFFFFFF; assign b = 64'h527FFFFFFFFFFFFF;

    #10 $display("\n2**728 * 2**295:");
    #10 assign a = 64'h6D70000000000000; assign b = 64'h5260000000000000;
    #10 assign a = 64'h6D7FFFFFFFFFFFFF; assign b = 64'h526FFFFFFFFFFFFF;

    #10 $display("\n2**729 * 2**294:");
    #10 assign a = 64'h6D80000000000000; assign b = 64'h5250000000000000;
    #10 assign a = 64'h6D8FFFFFFFFFFFFF; assign b = 64'h525FFFFFFFFFFFFF;

    #10 $display("\n2**730 * 2**293:");
    #10 assign a = 64'h6D90000000000000; assign b = 64'h5240000000000000;
    #10 assign a = 64'h6D9FFFFFFFFFFFFF; assign b = 64'h524FFFFFFFFFFFFF;

    #10 $display("\n2**731 * 2**292:");
    #10 assign a = 64'h6DA0000000000000; assign b = 64'h5230000000000000;
    #10 assign a = 64'h6DAFFFFFFFFFFFFF; assign b = 64'h523FFFFFFFFFFFFF;

    #10 $display("\n2**732 * 2**291:");
    #10 assign a = 64'h6DB0000000000000; assign b = 64'h5220000000000000;
    #10 assign a = 64'h6DBFFFFFFFFFFFFF; assign b = 64'h522FFFFFFFFFFFFF;

    #10 $display("\n2**733 * 2**290:");
    #10 assign a = 64'h6DC0000000000000; assign b = 64'h5210000000000000;
    #10 assign a = 64'h6DCFFFFFFFFFFFFF; assign b = 64'h521FFFFFFFFFFFFF;

    #10 $display("\n2**734 * 2**289:");
    #10 assign a = 64'h6DD0000000000000; assign b = 64'h5200000000000000;
    #10 assign a = 64'h6DDFFFFFFFFFFFFF; assign b = 64'h520FFFFFFFFFFFFF;

    #10 $display("\n2**735 * 2**288:");
    #10 assign a = 64'h6DE0000000000000; assign b = 64'h51F0000000000000;
    #10 assign a = 64'h6DEFFFFFFFFFFFFF; assign b = 64'h51FFFFFFFFFFFFFF;

    #10 $display("\n2**736 * 2**287:");
    #10 assign a = 64'h6DF0000000000000; assign b = 64'h51E0000000000000;
    #10 assign a = 64'h6DFFFFFFFFFFFFFF; assign b = 64'h51EFFFFFFFFFFFFF;

    #10 $display("\n2**737 * 2**286:");
    #10 assign a = 64'h6E00000000000000; assign b = 64'h51D0000000000000;
    #10 assign a = 64'h6E0FFFFFFFFFFFFF; assign b = 64'h51DFFFFFFFFFFFFF;

    #10 $display("\n2**738 * 2**285:");
    #10 assign a = 64'h6E10000000000000; assign b = 64'h51C0000000000000;
    #10 assign a = 64'h6E1FFFFFFFFFFFFF; assign b = 64'h51CFFFFFFFFFFFFF;

    #10 $display("\n2**739 * 2**284:");
    #10 assign a = 64'h6E20000000000000; assign b = 64'h51B0000000000000;
    #10 assign a = 64'h6E2FFFFFFFFFFFFF; assign b = 64'h51BFFFFFFFFFFFFF;

    #10 $display("\n2**740 * 2**283:");
    #10 assign a = 64'h6E30000000000000; assign b = 64'h51A0000000000000;
    #10 assign a = 64'h6E3FFFFFFFFFFFFF; assign b = 64'h51AFFFFFFFFFFFFF;

    #10 $display("\n2**741 * 2**282:");
    #10 assign a = 64'h6E40000000000000; assign b = 64'h5190000000000000;
    #10 assign a = 64'h6E4FFFFFFFFFFFFF; assign b = 64'h519FFFFFFFFFFFFF;

    #10 $display("\n2**742 * 2**281:");
    #10 assign a = 64'h6E50000000000000; assign b = 64'h5180000000000000;
    #10 assign a = 64'h6E5FFFFFFFFFFFFF; assign b = 64'h518FFFFFFFFFFFFF;

    #10 $display("\n2**743 * 2**280:");
    #10 assign a = 64'h6E60000000000000; assign b = 64'h5170000000000000;
    #10 assign a = 64'h6E6FFFFFFFFFFFFF; assign b = 64'h517FFFFFFFFFFFFF;

    #10 $display("\n2**744 * 2**279:");
    #10 assign a = 64'h6E70000000000000; assign b = 64'h5160000000000000;
    #10 assign a = 64'h6E7FFFFFFFFFFFFF; assign b = 64'h516FFFFFFFFFFFFF;

    #10 $display("\n2**745 * 2**278:");
    #10 assign a = 64'h6E80000000000000; assign b = 64'h5150000000000000;
    #10 assign a = 64'h6E8FFFFFFFFFFFFF; assign b = 64'h515FFFFFFFFFFFFF;

    #10 $display("\n2**746 * 2**277:");
    #10 assign a = 64'h6E90000000000000; assign b = 64'h5140000000000000;
    #10 assign a = 64'h6E9FFFFFFFFFFFFF; assign b = 64'h514FFFFFFFFFFFFF;

    #10 $display("\n2**747 * 2**276:");
    #10 assign a = 64'h6EA0000000000000; assign b = 64'h5130000000000000;
    #10 assign a = 64'h6EAFFFFFFFFFFFFF; assign b = 64'h513FFFFFFFFFFFFF;

    #10 $display("\n2**748 * 2**275:");
    #10 assign a = 64'h6EB0000000000000; assign b = 64'h5120000000000000;
    #10 assign a = 64'h6EBFFFFFFFFFFFFF; assign b = 64'h512FFFFFFFFFFFFF;

    #10 $display("\n2**749 * 2**274:");
    #10 assign a = 64'h6EC0000000000000; assign b = 64'h5110000000000000;
    #10 assign a = 64'h6ECFFFFFFFFFFFFF; assign b = 64'h511FFFFFFFFFFFFF;

    #10 $display("\n2**750 * 2**273:");
    #10 assign a = 64'h6ED0000000000000; assign b = 64'h5100000000000000;
    #10 assign a = 64'h6EDFFFFFFFFFFFFF; assign b = 64'h510FFFFFFFFFFFFF;

    #10 $display("\n2**751 * 2**272:");
    #10 assign a = 64'h6EE0000000000000; assign b = 64'h50F0000000000000;
    #10 assign a = 64'h6EEFFFFFFFFFFFFF; assign b = 64'h50FFFFFFFFFFFFFF;

    #10 $display("\n2**752 * 2**271:");
    #10 assign a = 64'h6EF0000000000000; assign b = 64'h50E0000000000000;
    #10 assign a = 64'h6EFFFFFFFFFFFFFF; assign b = 64'h50EFFFFFFFFFFFFF;

    #10 $display("\n2**753 * 2**270:");
    #10 assign a = 64'h6F00000000000000; assign b = 64'h50D0000000000000;
    #10 assign a = 64'h6F0FFFFFFFFFFFFF; assign b = 64'h50DFFFFFFFFFFFFF;

    #10 $display("\n2**754 * 2**269:");
    #10 assign a = 64'h6F10000000000000; assign b = 64'h50C0000000000000;
    #10 assign a = 64'h6F1FFFFFFFFFFFFF; assign b = 64'h50CFFFFFFFFFFFFF;

    #10 $display("\n2**755 * 2**268:");
    #10 assign a = 64'h6F20000000000000; assign b = 64'h50B0000000000000;
    #10 assign a = 64'h6F2FFFFFFFFFFFFF; assign b = 64'h50BFFFFFFFFFFFFF;

    #10 $display("\n2**756 * 2**267:");
    #10 assign a = 64'h6F30000000000000; assign b = 64'h50A0000000000000;
    #10 assign a = 64'h6F3FFFFFFFFFFFFF; assign b = 64'h50AFFFFFFFFFFFFF;

    #10 $display("\n2**757 * 2**266:");
    #10 assign a = 64'h6F40000000000000; assign b = 64'h5090000000000000;
    #10 assign a = 64'h6F4FFFFFFFFFFFFF; assign b = 64'h509FFFFFFFFFFFFF;

    #10 $display("\n2**758 * 2**265:");
    #10 assign a = 64'h6F50000000000000; assign b = 64'h5080000000000000;
    #10 assign a = 64'h6F5FFFFFFFFFFFFF; assign b = 64'h508FFFFFFFFFFFFF;

    #10 $display("\n2**759 * 2**264:");
    #10 assign a = 64'h6F60000000000000; assign b = 64'h5070000000000000;
    #10 assign a = 64'h6F6FFFFFFFFFFFFF; assign b = 64'h507FFFFFFFFFFFFF;

    #10 $display("\n2**760 * 2**263:");
    #10 assign a = 64'h6F70000000000000; assign b = 64'h5060000000000000;
    #10 assign a = 64'h6F7FFFFFFFFFFFFF; assign b = 64'h506FFFFFFFFFFFFF;

    #10 $display("\n2**761 * 2**262:");
    #10 assign a = 64'h6F80000000000000; assign b = 64'h5050000000000000;
    #10 assign a = 64'h6F8FFFFFFFFFFFFF; assign b = 64'h505FFFFFFFFFFFFF;

    #10 $display("\n2**762 * 2**261:");
    #10 assign a = 64'h6F90000000000000; assign b = 64'h5040000000000000;
    #10 assign a = 64'h6F9FFFFFFFFFFFFF; assign b = 64'h504FFFFFFFFFFFFF;

    #10 $display("\n2**763 * 2**260:");
    #10 assign a = 64'h6FA0000000000000; assign b = 64'h5030000000000000;
    #10 assign a = 64'h6FAFFFFFFFFFFFFF; assign b = 64'h503FFFFFFFFFFFFF;

    #10 $display("\n2**764 * 2**259:");
    #10 assign a = 64'h6FB0000000000000; assign b = 64'h5020000000000000;
    #10 assign a = 64'h6FBFFFFFFFFFFFFF; assign b = 64'h502FFFFFFFFFFFFF;

    #10 $display("\n2**765 * 2**258:");
    #10 assign a = 64'h6FC0000000000000; assign b = 64'h5010000000000000;
    #10 assign a = 64'h6FCFFFFFFFFFFFFF; assign b = 64'h501FFFFFFFFFFFFF;

    #10 $display("\n2**766 * 2**257:");
    #10 assign a = 64'h6FD0000000000000; assign b = 64'h5000000000000000;
    #10 assign a = 64'h6FDFFFFFFFFFFFFF; assign b = 64'h500FFFFFFFFFFFFF;

    #10 $display("\n2**767 * 2**256:");
    #10 assign a = 64'h6FE0000000000000; assign b = 64'h4FF0000000000000;
    #10 assign a = 64'h6FEFFFFFFFFFFFFF; assign b = 64'h4FFFFFFFFFFFFFFF;

    #10 $display("\n2**768 * 2**255:");
    #10 assign a = 64'h6FF0000000000000; assign b = 64'h4FE0000000000000;
    #10 assign a = 64'h6FFFFFFFFFFFFFFF; assign b = 64'h4FEFFFFFFFFFFFFF;

    #10 $display("\n2**769 * 2**254:");
    #10 assign a = 64'h7000000000000000; assign b = 64'h4FD0000000000000;
    #10 assign a = 64'h700FFFFFFFFFFFFF; assign b = 64'h4FDFFFFFFFFFFFFF;

    #10 $display("\n2**770 * 2**253:");
    #10 assign a = 64'h7010000000000000; assign b = 64'h4FC0000000000000;
    #10 assign a = 64'h701FFFFFFFFFFFFF; assign b = 64'h4FCFFFFFFFFFFFFF;

    #10 $display("\n2**771 * 2**252:");
    #10 assign a = 64'h7020000000000000; assign b = 64'h4FB0000000000000;
    #10 assign a = 64'h702FFFFFFFFFFFFF; assign b = 64'h4FBFFFFFFFFFFFFF;

    #10 $display("\n2**772 * 2**251:");
    #10 assign a = 64'h7030000000000000; assign b = 64'h4FA0000000000000;
    #10 assign a = 64'h703FFFFFFFFFFFFF; assign b = 64'h4FAFFFFFFFFFFFFF;

    #10 $display("\n2**773 * 2**250:");
    #10 assign a = 64'h7040000000000000; assign b = 64'h4F90000000000000;
    #10 assign a = 64'h704FFFFFFFFFFFFF; assign b = 64'h4F9FFFFFFFFFFFFF;

    #10 $display("\n2**774 * 2**249:");
    #10 assign a = 64'h7050000000000000; assign b = 64'h4F80000000000000;
    #10 assign a = 64'h705FFFFFFFFFFFFF; assign b = 64'h4F8FFFFFFFFFFFFF;

    #10 $display("\n2**775 * 2**248:");
    #10 assign a = 64'h7060000000000000; assign b = 64'h4F70000000000000;
    #10 assign a = 64'h706FFFFFFFFFFFFF; assign b = 64'h4F7FFFFFFFFFFFFF;

    #10 $display("\n2**776 * 2**247:");
    #10 assign a = 64'h7070000000000000; assign b = 64'h4F60000000000000;
    #10 assign a = 64'h707FFFFFFFFFFFFF; assign b = 64'h4F6FFFFFFFFFFFFF;

    #10 $display("\n2**777 * 2**246:");
    #10 assign a = 64'h7080000000000000; assign b = 64'h4F50000000000000;
    #10 assign a = 64'h708FFFFFFFFFFFFF; assign b = 64'h4F5FFFFFFFFFFFFF;

    #10 $display("\n2**778 * 2**245:");
    #10 assign a = 64'h7090000000000000; assign b = 64'h4F40000000000000;
    #10 assign a = 64'h709FFFFFFFFFFFFF; assign b = 64'h4F4FFFFFFFFFFFFF;

    #10 $display("\n2**779 * 2**244:");
    #10 assign a = 64'h70A0000000000000; assign b = 64'h4F30000000000000;
    #10 assign a = 64'h70AFFFFFFFFFFFFF; assign b = 64'h4F3FFFFFFFFFFFFF;

    #10 $display("\n2**780 * 2**243:");
    #10 assign a = 64'h70B0000000000000; assign b = 64'h4F20000000000000;
    #10 assign a = 64'h70BFFFFFFFFFFFFF; assign b = 64'h4F2FFFFFFFFFFFFF;

    #10 $display("\n2**781 * 2**242:");
    #10 assign a = 64'h70C0000000000000; assign b = 64'h4F10000000000000;
    #10 assign a = 64'h70CFFFFFFFFFFFFF; assign b = 64'h4F1FFFFFFFFFFFFF;

    #10 $display("\n2**782 * 2**241:");
    #10 assign a = 64'h70D0000000000000; assign b = 64'h4F00000000000000;
    #10 assign a = 64'h70DFFFFFFFFFFFFF; assign b = 64'h4F0FFFFFFFFFFFFF;

    #10 $display("\n2**783 * 2**240:");
    #10 assign a = 64'h70E0000000000000; assign b = 64'h4EF0000000000000;
    #10 assign a = 64'h70EFFFFFFFFFFFFF; assign b = 64'h4EFFFFFFFFFFFFFF;

    #10 $display("\n2**784 * 2**239:");
    #10 assign a = 64'h70F0000000000000; assign b = 64'h4EE0000000000000;
    #10 assign a = 64'h70FFFFFFFFFFFFFF; assign b = 64'h4EEFFFFFFFFFFFFF;

    #10 $display("\n2**785 * 2**238:");
    #10 assign a = 64'h7100000000000000; assign b = 64'h4ED0000000000000;
    #10 assign a = 64'h710FFFFFFFFFFFFF; assign b = 64'h4EDFFFFFFFFFFFFF;

    #10 $display("\n2**786 * 2**237:");
    #10 assign a = 64'h7110000000000000; assign b = 64'h4EC0000000000000;
    #10 assign a = 64'h711FFFFFFFFFFFFF; assign b = 64'h4ECFFFFFFFFFFFFF;

    #10 $display("\n2**787 * 2**236:");
    #10 assign a = 64'h7120000000000000; assign b = 64'h4EB0000000000000;
    #10 assign a = 64'h712FFFFFFFFFFFFF; assign b = 64'h4EBFFFFFFFFFFFFF;

    #10 $display("\n2**788 * 2**235:");
    #10 assign a = 64'h7130000000000000; assign b = 64'h4EA0000000000000;
    #10 assign a = 64'h713FFFFFFFFFFFFF; assign b = 64'h4EAFFFFFFFFFFFFF;

    #10 $display("\n2**789 * 2**234:");
    #10 assign a = 64'h7140000000000000; assign b = 64'h4E90000000000000;
    #10 assign a = 64'h714FFFFFFFFFFFFF; assign b = 64'h4E9FFFFFFFFFFFFF;

    #10 $display("\n2**790 * 2**233:");
    #10 assign a = 64'h7150000000000000; assign b = 64'h4E80000000000000;
    #10 assign a = 64'h715FFFFFFFFFFFFF; assign b = 64'h4E8FFFFFFFFFFFFF;

    #10 $display("\n2**791 * 2**232:");
    #10 assign a = 64'h7160000000000000; assign b = 64'h4E70000000000000;
    #10 assign a = 64'h716FFFFFFFFFFFFF; assign b = 64'h4E7FFFFFFFFFFFFF;

    #10 $display("\n2**792 * 2**231:");
    #10 assign a = 64'h7170000000000000; assign b = 64'h4E60000000000000;
    #10 assign a = 64'h717FFFFFFFFFFFFF; assign b = 64'h4E6FFFFFFFFFFFFF;

    #10 $display("\n2**793 * 2**230:");
    #10 assign a = 64'h7180000000000000; assign b = 64'h4E50000000000000;
    #10 assign a = 64'h718FFFFFFFFFFFFF; assign b = 64'h4E5FFFFFFFFFFFFF;

    #10 $display("\n2**794 * 2**229:");
    #10 assign a = 64'h7190000000000000; assign b = 64'h4E40000000000000;
    #10 assign a = 64'h719FFFFFFFFFFFFF; assign b = 64'h4E4FFFFFFFFFFFFF;

    #10 $display("\n2**795 * 2**228:");
    #10 assign a = 64'h71A0000000000000; assign b = 64'h4E30000000000000;
    #10 assign a = 64'h71AFFFFFFFFFFFFF; assign b = 64'h4E3FFFFFFFFFFFFF;

    #10 $display("\n2**796 * 2**227:");
    #10 assign a = 64'h71B0000000000000; assign b = 64'h4E20000000000000;
    #10 assign a = 64'h71BFFFFFFFFFFFFF; assign b = 64'h4E2FFFFFFFFFFFFF;

    #10 $display("\n2**797 * 2**226:");
    #10 assign a = 64'h71C0000000000000; assign b = 64'h4E10000000000000;
    #10 assign a = 64'h71CFFFFFFFFFFFFF; assign b = 64'h4E1FFFFFFFFFFFFF;

    #10 $display("\n2**798 * 2**225:");
    #10 assign a = 64'h71D0000000000000; assign b = 64'h4E00000000000000;
    #10 assign a = 64'h71DFFFFFFFFFFFFF; assign b = 64'h4E0FFFFFFFFFFFFF;

    #10 $display("\n2**799 * 2**224:");
    #10 assign a = 64'h71E0000000000000; assign b = 64'h4DF0000000000000;
    #10 assign a = 64'h71EFFFFFFFFFFFFF; assign b = 64'h4DFFFFFFFFFFFFFF;

    #10 $display("\n2**800 * 2**223:");
    #10 assign a = 64'h71F0000000000000; assign b = 64'h4DE0000000000000;
    #10 assign a = 64'h71FFFFFFFFFFFFFF; assign b = 64'h4DEFFFFFFFFFFFFF;

    #10 $display("\n2**801 * 2**222:");
    #10 assign a = 64'h7200000000000000; assign b = 64'h4DD0000000000000;
    #10 assign a = 64'h720FFFFFFFFFFFFF; assign b = 64'h4DDFFFFFFFFFFFFF;

    #10 $display("\n2**802 * 2**221:");
    #10 assign a = 64'h7210000000000000; assign b = 64'h4DC0000000000000;
    #10 assign a = 64'h721FFFFFFFFFFFFF; assign b = 64'h4DCFFFFFFFFFFFFF;

    #10 $display("\n2**803 * 2**220:");
    #10 assign a = 64'h7220000000000000; assign b = 64'h4DB0000000000000;
    #10 assign a = 64'h722FFFFFFFFFFFFF; assign b = 64'h4DBFFFFFFFFFFFFF;

    #10 $display("\n2**804 * 2**219:");
    #10 assign a = 64'h7230000000000000; assign b = 64'h4DA0000000000000;
    #10 assign a = 64'h723FFFFFFFFFFFFF; assign b = 64'h4DAFFFFFFFFFFFFF;

    #10 $display("\n2**805 * 2**218:");
    #10 assign a = 64'h7240000000000000; assign b = 64'h4D90000000000000;
    #10 assign a = 64'h724FFFFFFFFFFFFF; assign b = 64'h4D9FFFFFFFFFFFFF;

    #10 $display("\n2**806 * 2**217:");
    #10 assign a = 64'h7250000000000000; assign b = 64'h4D80000000000000;
    #10 assign a = 64'h725FFFFFFFFFFFFF; assign b = 64'h4D8FFFFFFFFFFFFF;

    #10 $display("\n2**807 * 2**216:");
    #10 assign a = 64'h7260000000000000; assign b = 64'h4D70000000000000;
    #10 assign a = 64'h726FFFFFFFFFFFFF; assign b = 64'h4D7FFFFFFFFFFFFF;

    #10 $display("\n2**808 * 2**215:");
    #10 assign a = 64'h7270000000000000; assign b = 64'h4D60000000000000;
    #10 assign a = 64'h727FFFFFFFFFFFFF; assign b = 64'h4D6FFFFFFFFFFFFF;

    #10 $display("\n2**809 * 2**214:");
    #10 assign a = 64'h7280000000000000; assign b = 64'h4D50000000000000;
    #10 assign a = 64'h728FFFFFFFFFFFFF; assign b = 64'h4D5FFFFFFFFFFFFF;

    #10 $display("\n2**810 * 2**213:");
    #10 assign a = 64'h7290000000000000; assign b = 64'h4D40000000000000;
    #10 assign a = 64'h729FFFFFFFFFFFFF; assign b = 64'h4D4FFFFFFFFFFFFF;

    #10 $display("\n2**811 * 2**212:");
    #10 assign a = 64'h72A0000000000000; assign b = 64'h4D30000000000000;
    #10 assign a = 64'h72AFFFFFFFFFFFFF; assign b = 64'h4D3FFFFFFFFFFFFF;

    #10 $display("\n2**812 * 2**211:");
    #10 assign a = 64'h72B0000000000000; assign b = 64'h4D20000000000000;
    #10 assign a = 64'h72BFFFFFFFFFFFFF; assign b = 64'h4D2FFFFFFFFFFFFF;

    #10 $display("\n2**813 * 2**210:");
    #10 assign a = 64'h72C0000000000000; assign b = 64'h4D10000000000000;
    #10 assign a = 64'h72CFFFFFFFFFFFFF; assign b = 64'h4D1FFFFFFFFFFFFF;

    #10 $display("\n2**814 * 2**209:");
    #10 assign a = 64'h72D0000000000000; assign b = 64'h4D00000000000000;
    #10 assign a = 64'h72DFFFFFFFFFFFFF; assign b = 64'h4D0FFFFFFFFFFFFF;

    #10 $display("\n2**815 * 2**208:");
    #10 assign a = 64'h72E0000000000000; assign b = 64'h4CF0000000000000;
    #10 assign a = 64'h72EFFFFFFFFFFFFF; assign b = 64'h4CFFFFFFFFFFFFFF;

    #10 $display("\n2**816 * 2**207:");
    #10 assign a = 64'h72F0000000000000; assign b = 64'h4CE0000000000000;
    #10 assign a = 64'h72FFFFFFFFFFFFFF; assign b = 64'h4CEFFFFFFFFFFFFF;

    #10 $display("\n2**817 * 2**206:");
    #10 assign a = 64'h7300000000000000; assign b = 64'h4CD0000000000000;
    #10 assign a = 64'h730FFFFFFFFFFFFF; assign b = 64'h4CDFFFFFFFFFFFFF;

    #10 $display("\n2**818 * 2**205:");
    #10 assign a = 64'h7310000000000000; assign b = 64'h4CC0000000000000;
    #10 assign a = 64'h731FFFFFFFFFFFFF; assign b = 64'h4CCFFFFFFFFFFFFF;

    #10 $display("\n2**819 * 2**204:");
    #10 assign a = 64'h7320000000000000; assign b = 64'h4CB0000000000000;
    #10 assign a = 64'h732FFFFFFFFFFFFF; assign b = 64'h4CBFFFFFFFFFFFFF;

    #10 $display("\n2**820 * 2**203:");
    #10 assign a = 64'h7330000000000000; assign b = 64'h4CA0000000000000;
    #10 assign a = 64'h733FFFFFFFFFFFFF; assign b = 64'h4CAFFFFFFFFFFFFF;

    #10 $display("\n2**821 * 2**202:");
    #10 assign a = 64'h7340000000000000; assign b = 64'h4C90000000000000;
    #10 assign a = 64'h734FFFFFFFFFFFFF; assign b = 64'h4C9FFFFFFFFFFFFF;

    #10 $display("\n2**822 * 2**201:");
    #10 assign a = 64'h7350000000000000; assign b = 64'h4C80000000000000;
    #10 assign a = 64'h735FFFFFFFFFFFFF; assign b = 64'h4C8FFFFFFFFFFFFF;

    #10 $display("\n2**823 * 2**200:");
    #10 assign a = 64'h7360000000000000; assign b = 64'h4C70000000000000;
    #10 assign a = 64'h736FFFFFFFFFFFFF; assign b = 64'h4C7FFFFFFFFFFFFF;

    #10 $display("\n2**824 * 2**199:");
    #10 assign a = 64'h7370000000000000; assign b = 64'h4C60000000000000;
    #10 assign a = 64'h737FFFFFFFFFFFFF; assign b = 64'h4C6FFFFFFFFFFFFF;

    #10 $display("\n2**825 * 2**198:");
    #10 assign a = 64'h7380000000000000; assign b = 64'h4C50000000000000;
    #10 assign a = 64'h738FFFFFFFFFFFFF; assign b = 64'h4C5FFFFFFFFFFFFF;

    #10 $display("\n2**826 * 2**197:");
    #10 assign a = 64'h7390000000000000; assign b = 64'h4C40000000000000;
    #10 assign a = 64'h739FFFFFFFFFFFFF; assign b = 64'h4C4FFFFFFFFFFFFF;

    #10 $display("\n2**827 * 2**196:");
    #10 assign a = 64'h73A0000000000000; assign b = 64'h4C30000000000000;
    #10 assign a = 64'h73AFFFFFFFFFFFFF; assign b = 64'h4C3FFFFFFFFFFFFF;

    #10 $display("\n2**828 * 2**195:");
    #10 assign a = 64'h73B0000000000000; assign b = 64'h4C20000000000000;
    #10 assign a = 64'h73BFFFFFFFFFFFFF; assign b = 64'h4C2FFFFFFFFFFFFF;

    #10 $display("\n2**829 * 2**194:");
    #10 assign a = 64'h73C0000000000000; assign b = 64'h4C10000000000000;
    #10 assign a = 64'h73CFFFFFFFFFFFFF; assign b = 64'h4C1FFFFFFFFFFFFF;

    #10 $display("\n2**830 * 2**193:");
    #10 assign a = 64'h73D0000000000000; assign b = 64'h4C00000000000000;
    #10 assign a = 64'h73DFFFFFFFFFFFFF; assign b = 64'h4C0FFFFFFFFFFFFF;

    #10 $display("\n2**831 * 2**192:");
    #10 assign a = 64'h73E0000000000000; assign b = 64'h4BF0000000000000;
    #10 assign a = 64'h73EFFFFFFFFFFFFF; assign b = 64'h4BFFFFFFFFFFFFFF;

    #10 $display("\n2**832 * 2**191:");
    #10 assign a = 64'h73F0000000000000; assign b = 64'h4BE0000000000000;
    #10 assign a = 64'h73FFFFFFFFFFFFFF; assign b = 64'h4BEFFFFFFFFFFFFF;

    #10 $display("\n2**833 * 2**190:");
    #10 assign a = 64'h7400000000000000; assign b = 64'h4BD0000000000000;
    #10 assign a = 64'h740FFFFFFFFFFFFF; assign b = 64'h4BDFFFFFFFFFFFFF;

    #10 $display("\n2**834 * 2**189:");
    #10 assign a = 64'h7410000000000000; assign b = 64'h4BC0000000000000;
    #10 assign a = 64'h741FFFFFFFFFFFFF; assign b = 64'h4BCFFFFFFFFFFFFF;

    #10 $display("\n2**835 * 2**188:");
    #10 assign a = 64'h7420000000000000; assign b = 64'h4BB0000000000000;
    #10 assign a = 64'h742FFFFFFFFFFFFF; assign b = 64'h4BBFFFFFFFFFFFFF;

    #10 $display("\n2**836 * 2**187:");
    #10 assign a = 64'h7430000000000000; assign b = 64'h4BA0000000000000;
    #10 assign a = 64'h743FFFFFFFFFFFFF; assign b = 64'h4BAFFFFFFFFFFFFF;

    #10 $display("\n2**837 * 2**186:");
    #10 assign a = 64'h7440000000000000; assign b = 64'h4B90000000000000;
    #10 assign a = 64'h744FFFFFFFFFFFFF; assign b = 64'h4B9FFFFFFFFFFFFF;

    #10 $display("\n2**838 * 2**185:");
    #10 assign a = 64'h7450000000000000; assign b = 64'h4B80000000000000;
    #10 assign a = 64'h745FFFFFFFFFFFFF; assign b = 64'h4B8FFFFFFFFFFFFF;

    #10 $display("\n2**839 * 2**184:");
    #10 assign a = 64'h7460000000000000; assign b = 64'h4B70000000000000;
    #10 assign a = 64'h746FFFFFFFFFFFFF; assign b = 64'h4B7FFFFFFFFFFFFF;

    #10 $display("\n2**840 * 2**183:");
    #10 assign a = 64'h7470000000000000; assign b = 64'h4B60000000000000;
    #10 assign a = 64'h747FFFFFFFFFFFFF; assign b = 64'h4B6FFFFFFFFFFFFF;

    #10 $display("\n2**841 * 2**182:");
    #10 assign a = 64'h7480000000000000; assign b = 64'h4B50000000000000;
    #10 assign a = 64'h748FFFFFFFFFFFFF; assign b = 64'h4B5FFFFFFFFFFFFF;

    #10 $display("\n2**842 * 2**181:");
    #10 assign a = 64'h7490000000000000; assign b = 64'h4B40000000000000;
    #10 assign a = 64'h749FFFFFFFFFFFFF; assign b = 64'h4B4FFFFFFFFFFFFF;

    #10 $display("\n2**843 * 2**180:");
    #10 assign a = 64'h74A0000000000000; assign b = 64'h4B30000000000000;
    #10 assign a = 64'h74AFFFFFFFFFFFFF; assign b = 64'h4B3FFFFFFFFFFFFF;

    #10 $display("\n2**844 * 2**179:");
    #10 assign a = 64'h74B0000000000000; assign b = 64'h4B20000000000000;
    #10 assign a = 64'h74BFFFFFFFFFFFFF; assign b = 64'h4B2FFFFFFFFFFFFF;

    #10 $display("\n2**845 * 2**178:");
    #10 assign a = 64'h74C0000000000000; assign b = 64'h4B10000000000000;
    #10 assign a = 64'h74CFFFFFFFFFFFFF; assign b = 64'h4B1FFFFFFFFFFFFF;

    #10 $display("\n2**846 * 2**177:");
    #10 assign a = 64'h74D0000000000000; assign b = 64'h4B00000000000000;
    #10 assign a = 64'h74DFFFFFFFFFFFFF; assign b = 64'h4B0FFFFFFFFFFFFF;

    #10 $display("\n2**847 * 2**176:");
    #10 assign a = 64'h74E0000000000000; assign b = 64'h4AF0000000000000;
    #10 assign a = 64'h74EFFFFFFFFFFFFF; assign b = 64'h4AFFFFFFFFFFFFFF;

    #10 $display("\n2**848 * 2**175:");
    #10 assign a = 64'h74F0000000000000; assign b = 64'h4AE0000000000000;
    #10 assign a = 64'h74FFFFFFFFFFFFFF; assign b = 64'h4AEFFFFFFFFFFFFF;

    #10 $display("\n2**849 * 2**174:");
    #10 assign a = 64'h7500000000000000; assign b = 64'h4AD0000000000000;
    #10 assign a = 64'h750FFFFFFFFFFFFF; assign b = 64'h4ADFFFFFFFFFFFFF;

    #10 $display("\n2**850 * 2**173:");
    #10 assign a = 64'h7510000000000000; assign b = 64'h4AC0000000000000;
    #10 assign a = 64'h751FFFFFFFFFFFFF; assign b = 64'h4ACFFFFFFFFFFFFF;

    #10 $display("\n2**851 * 2**172:");
    #10 assign a = 64'h7520000000000000; assign b = 64'h4AB0000000000000;
    #10 assign a = 64'h752FFFFFFFFFFFFF; assign b = 64'h4ABFFFFFFFFFFFFF;

    #10 $display("\n2**852 * 2**171:");
    #10 assign a = 64'h7530000000000000; assign b = 64'h4AA0000000000000;
    #10 assign a = 64'h753FFFFFFFFFFFFF; assign b = 64'h4AAFFFFFFFFFFFFF;

    #10 $display("\n2**853 * 2**170:");
    #10 assign a = 64'h7540000000000000; assign b = 64'h4A90000000000000;
    #10 assign a = 64'h754FFFFFFFFFFFFF; assign b = 64'h4A9FFFFFFFFFFFFF;

    #10 $display("\n2**854 * 2**169:");
    #10 assign a = 64'h7550000000000000; assign b = 64'h4A80000000000000;
    #10 assign a = 64'h755FFFFFFFFFFFFF; assign b = 64'h4A8FFFFFFFFFFFFF;

    #10 $display("\n2**855 * 2**168:");
    #10 assign a = 64'h7560000000000000; assign b = 64'h4A70000000000000;
    #10 assign a = 64'h756FFFFFFFFFFFFF; assign b = 64'h4A7FFFFFFFFFFFFF;

    #10 $display("\n2**856 * 2**167:");
    #10 assign a = 64'h7570000000000000; assign b = 64'h4A60000000000000;
    #10 assign a = 64'h757FFFFFFFFFFFFF; assign b = 64'h4A6FFFFFFFFFFFFF;

    #10 $display("\n2**857 * 2**166:");
    #10 assign a = 64'h7580000000000000; assign b = 64'h4A50000000000000;
    #10 assign a = 64'h758FFFFFFFFFFFFF; assign b = 64'h4A5FFFFFFFFFFFFF;

    #10 $display("\n2**858 * 2**165:");
    #10 assign a = 64'h7590000000000000; assign b = 64'h4A40000000000000;
    #10 assign a = 64'h759FFFFFFFFFFFFF; assign b = 64'h4A4FFFFFFFFFFFFF;

    #10 $display("\n2**859 * 2**164:");
    #10 assign a = 64'h75A0000000000000; assign b = 64'h4A30000000000000;
    #10 assign a = 64'h75AFFFFFFFFFFFFF; assign b = 64'h4A3FFFFFFFFFFFFF;

    #10 $display("\n2**860 * 2**163:");
    #10 assign a = 64'h75B0000000000000; assign b = 64'h4A20000000000000;
    #10 assign a = 64'h75BFFFFFFFFFFFFF; assign b = 64'h4A2FFFFFFFFFFFFF;

    #10 $display("\n2**861 * 2**162:");
    #10 assign a = 64'h75C0000000000000; assign b = 64'h4A10000000000000;
    #10 assign a = 64'h75CFFFFFFFFFFFFF; assign b = 64'h4A1FFFFFFFFFFFFF;

    #10 $display("\n2**862 * 2**161:");
    #10 assign a = 64'h75D0000000000000; assign b = 64'h4A00000000000000;
    #10 assign a = 64'h75DFFFFFFFFFFFFF; assign b = 64'h4A0FFFFFFFFFFFFF;

    #10 $display("\n2**863 * 2**160:");
    #10 assign a = 64'h75E0000000000000; assign b = 64'h49F0000000000000;
    #10 assign a = 64'h75EFFFFFFFFFFFFF; assign b = 64'h49FFFFFFFFFFFFFF;

    #10 $display("\n2**864 * 2**159:");
    #10 assign a = 64'h75F0000000000000; assign b = 64'h49E0000000000000;
    #10 assign a = 64'h75FFFFFFFFFFFFFF; assign b = 64'h49EFFFFFFFFFFFFF;

    #10 $display("\n2**865 * 2**158:");
    #10 assign a = 64'h7600000000000000; assign b = 64'h49D0000000000000;
    #10 assign a = 64'h760FFFFFFFFFFFFF; assign b = 64'h49DFFFFFFFFFFFFF;

    #10 $display("\n2**866 * 2**157:");
    #10 assign a = 64'h7610000000000000; assign b = 64'h49C0000000000000;
    #10 assign a = 64'h761FFFFFFFFFFFFF; assign b = 64'h49CFFFFFFFFFFFFF;

    #10 $display("\n2**867 * 2**156:");
    #10 assign a = 64'h7620000000000000; assign b = 64'h49B0000000000000;
    #10 assign a = 64'h762FFFFFFFFFFFFF; assign b = 64'h49BFFFFFFFFFFFFF;

    #10 $display("\n2**868 * 2**155:");
    #10 assign a = 64'h7630000000000000; assign b = 64'h49A0000000000000;
    #10 assign a = 64'h763FFFFFFFFFFFFF; assign b = 64'h49AFFFFFFFFFFFFF;

    #10 $display("\n2**869 * 2**154:");
    #10 assign a = 64'h7640000000000000; assign b = 64'h4990000000000000;
    #10 assign a = 64'h764FFFFFFFFFFFFF; assign b = 64'h499FFFFFFFFFFFFF;

    #10 $display("\n2**870 * 2**153:");
    #10 assign a = 64'h7650000000000000; assign b = 64'h4980000000000000;
    #10 assign a = 64'h765FFFFFFFFFFFFF; assign b = 64'h498FFFFFFFFFFFFF;

    #10 $display("\n2**871 * 2**152:");
    #10 assign a = 64'h7660000000000000; assign b = 64'h4970000000000000;
    #10 assign a = 64'h766FFFFFFFFFFFFF; assign b = 64'h497FFFFFFFFFFFFF;

    #10 $display("\n2**872 * 2**151:");
    #10 assign a = 64'h7670000000000000; assign b = 64'h4960000000000000;
    #10 assign a = 64'h767FFFFFFFFFFFFF; assign b = 64'h496FFFFFFFFFFFFF;

    #10 $display("\n2**873 * 2**150:");
    #10 assign a = 64'h7680000000000000; assign b = 64'h4950000000000000;
    #10 assign a = 64'h768FFFFFFFFFFFFF; assign b = 64'h495FFFFFFFFFFFFF;

    #10 $display("\n2**874 * 2**149:");
    #10 assign a = 64'h7690000000000000; assign b = 64'h4940000000000000;
    #10 assign a = 64'h769FFFFFFFFFFFFF; assign b = 64'h494FFFFFFFFFFFFF;

    #10 $display("\n2**875 * 2**148:");
    #10 assign a = 64'h76A0000000000000; assign b = 64'h4930000000000000;
    #10 assign a = 64'h76AFFFFFFFFFFFFF; assign b = 64'h493FFFFFFFFFFFFF;

    #10 $display("\n2**876 * 2**147:");
    #10 assign a = 64'h76B0000000000000; assign b = 64'h4920000000000000;
    #10 assign a = 64'h76BFFFFFFFFFFFFF; assign b = 64'h492FFFFFFFFFFFFF;

    #10 $display("\n2**877 * 2**146:");
    #10 assign a = 64'h76C0000000000000; assign b = 64'h4910000000000000;
    #10 assign a = 64'h76CFFFFFFFFFFFFF; assign b = 64'h491FFFFFFFFFFFFF;

    #10 $display("\n2**878 * 2**145:");
    #10 assign a = 64'h76D0000000000000; assign b = 64'h4900000000000000;
    #10 assign a = 64'h76DFFFFFFFFFFFFF; assign b = 64'h490FFFFFFFFFFFFF;

    #10 $display("\n2**879 * 2**144:");
    #10 assign a = 64'h76E0000000000000; assign b = 64'h48F0000000000000;
    #10 assign a = 64'h76EFFFFFFFFFFFFF; assign b = 64'h48FFFFFFFFFFFFFF;

    #10 $display("\n2**880 * 2**143:");
    #10 assign a = 64'h76F0000000000000; assign b = 64'h48E0000000000000;
    #10 assign a = 64'h76FFFFFFFFFFFFFF; assign b = 64'h48EFFFFFFFFFFFFF;

    #10 $display("\n2**881 * 2**142:");
    #10 assign a = 64'h7700000000000000; assign b = 64'h48D0000000000000;
    #10 assign a = 64'h770FFFFFFFFFFFFF; assign b = 64'h48DFFFFFFFFFFFFF;

    #10 $display("\n2**882 * 2**141:");
    #10 assign a = 64'h7710000000000000; assign b = 64'h48C0000000000000;
    #10 assign a = 64'h771FFFFFFFFFFFFF; assign b = 64'h48CFFFFFFFFFFFFF;

    #10 $display("\n2**883 * 2**140:");
    #10 assign a = 64'h7720000000000000; assign b = 64'h48B0000000000000;
    #10 assign a = 64'h772FFFFFFFFFFFFF; assign b = 64'h48BFFFFFFFFFFFFF;

    #10 $display("\n2**884 * 2**139:");
    #10 assign a = 64'h7730000000000000; assign b = 64'h48A0000000000000;
    #10 assign a = 64'h773FFFFFFFFFFFFF; assign b = 64'h48AFFFFFFFFFFFFF;

    #10 $display("\n2**885 * 2**138:");
    #10 assign a = 64'h7740000000000000; assign b = 64'h4890000000000000;
    #10 assign a = 64'h774FFFFFFFFFFFFF; assign b = 64'h489FFFFFFFFFFFFF;

    #10 $display("\n2**886 * 2**137:");
    #10 assign a = 64'h7750000000000000; assign b = 64'h4880000000000000;
    #10 assign a = 64'h775FFFFFFFFFFFFF; assign b = 64'h488FFFFFFFFFFFFF;

    #10 $display("\n2**887 * 2**136:");
    #10 assign a = 64'h7760000000000000; assign b = 64'h4870000000000000;
    #10 assign a = 64'h776FFFFFFFFFFFFF; assign b = 64'h487FFFFFFFFFFFFF;

    #10 $display("\n2**888 * 2**135:");
    #10 assign a = 64'h7770000000000000; assign b = 64'h4860000000000000;
    #10 assign a = 64'h777FFFFFFFFFFFFF; assign b = 64'h486FFFFFFFFFFFFF;

    #10 $display("\n2**889 * 2**134:");
    #10 assign a = 64'h7780000000000000; assign b = 64'h4850000000000000;
    #10 assign a = 64'h778FFFFFFFFFFFFF; assign b = 64'h485FFFFFFFFFFFFF;

    #10 $display("\n2**890 * 2**133:");
    #10 assign a = 64'h7790000000000000; assign b = 64'h4840000000000000;
    #10 assign a = 64'h779FFFFFFFFFFFFF; assign b = 64'h484FFFFFFFFFFFFF;

    #10 $display("\n2**891 * 2**132:");
    #10 assign a = 64'h77A0000000000000; assign b = 64'h4830000000000000;
    #10 assign a = 64'h77AFFFFFFFFFFFFF; assign b = 64'h483FFFFFFFFFFFFF;

    #10 $display("\n2**892 * 2**131:");
    #10 assign a = 64'h77B0000000000000; assign b = 64'h4820000000000000;
    #10 assign a = 64'h77BFFFFFFFFFFFFF; assign b = 64'h482FFFFFFFFFFFFF;

    #10 $display("\n2**893 * 2**130:");
    #10 assign a = 64'h77C0000000000000; assign b = 64'h4810000000000000;
    #10 assign a = 64'h77CFFFFFFFFFFFFF; assign b = 64'h481FFFFFFFFFFFFF;

    #10 $display("\n2**894 * 2**129:");
    #10 assign a = 64'h77D0000000000000; assign b = 64'h4800000000000000;
    #10 assign a = 64'h77DFFFFFFFFFFFFF; assign b = 64'h480FFFFFFFFFFFFF;

    #10 $display("\n2**895 * 2**128:");
    #10 assign a = 64'h77E0000000000000; assign b = 64'h47F0000000000000;
    #10 assign a = 64'h77EFFFFFFFFFFFFF; assign b = 64'h47FFFFFFFFFFFFFF;

    #10 $display("\n2**896 * 2**127:");
    #10 assign a = 64'h77F0000000000000; assign b = 64'h47E0000000000000;
    #10 assign a = 64'h77FFFFFFFFFFFFFF; assign b = 64'h47EFFFFFFFFFFFFF;

    #10 $display("\n2**897 * 2**126:");
    #10 assign a = 64'h7800000000000000; assign b = 64'h47D0000000000000;
    #10 assign a = 64'h780FFFFFFFFFFFFF; assign b = 64'h47DFFFFFFFFFFFFF;

    #10 $display("\n2**898 * 2**125:");
    #10 assign a = 64'h7810000000000000; assign b = 64'h47C0000000000000;
    #10 assign a = 64'h781FFFFFFFFFFFFF; assign b = 64'h47CFFFFFFFFFFFFF;

    #10 $display("\n2**899 * 2**124:");
    #10 assign a = 64'h7820000000000000; assign b = 64'h47B0000000000000;
    #10 assign a = 64'h782FFFFFFFFFFFFF; assign b = 64'h47BFFFFFFFFFFFFF;

    #10 $display("\n2**900 * 2**123:");
    #10 assign a = 64'h7830000000000000; assign b = 64'h47A0000000000000;
    #10 assign a = 64'h783FFFFFFFFFFFFF; assign b = 64'h47AFFFFFFFFFFFFF;

    #10 $display("\n2**901 * 2**122:");
    #10 assign a = 64'h7840000000000000; assign b = 64'h4790000000000000;
    #10 assign a = 64'h784FFFFFFFFFFFFF; assign b = 64'h479FFFFFFFFFFFFF;

    #10 $display("\n2**902 * 2**121:");
    #10 assign a = 64'h7850000000000000; assign b = 64'h4780000000000000;
    #10 assign a = 64'h785FFFFFFFFFFFFF; assign b = 64'h478FFFFFFFFFFFFF;

    #10 $display("\n2**903 * 2**120:");
    #10 assign a = 64'h7860000000000000; assign b = 64'h4770000000000000;
    #10 assign a = 64'h786FFFFFFFFFFFFF; assign b = 64'h477FFFFFFFFFFFFF;

    #10 $display("\n2**904 * 2**119:");
    #10 assign a = 64'h7870000000000000; assign b = 64'h4760000000000000;
    #10 assign a = 64'h787FFFFFFFFFFFFF; assign b = 64'h476FFFFFFFFFFFFF;

    #10 $display("\n2**905 * 2**118:");
    #10 assign a = 64'h7880000000000000; assign b = 64'h4750000000000000;
    #10 assign a = 64'h788FFFFFFFFFFFFF; assign b = 64'h475FFFFFFFFFFFFF;

    #10 $display("\n2**906 * 2**117:");
    #10 assign a = 64'h7890000000000000; assign b = 64'h4740000000000000;
    #10 assign a = 64'h789FFFFFFFFFFFFF; assign b = 64'h474FFFFFFFFFFFFF;

    #10 $display("\n2**907 * 2**116:");
    #10 assign a = 64'h78A0000000000000; assign b = 64'h4730000000000000;
    #10 assign a = 64'h78AFFFFFFFFFFFFF; assign b = 64'h473FFFFFFFFFFFFF;

    #10 $display("\n2**908 * 2**115:");
    #10 assign a = 64'h78B0000000000000; assign b = 64'h4720000000000000;
    #10 assign a = 64'h78BFFFFFFFFFFFFF; assign b = 64'h472FFFFFFFFFFFFF;

    #10 $display("\n2**909 * 2**114:");
    #10 assign a = 64'h78C0000000000000; assign b = 64'h4710000000000000;
    #10 assign a = 64'h78CFFFFFFFFFFFFF; assign b = 64'h471FFFFFFFFFFFFF;

    #10 $display("\n2**910 * 2**113:");
    #10 assign a = 64'h78D0000000000000; assign b = 64'h4700000000000000;
    #10 assign a = 64'h78DFFFFFFFFFFFFF; assign b = 64'h470FFFFFFFFFFFFF;

    #10 $display("\n2**911 * 2**112:");
    #10 assign a = 64'h78E0000000000000; assign b = 64'h46F0000000000000;
    #10 assign a = 64'h78EFFFFFFFFFFFFF; assign b = 64'h46FFFFFFFFFFFFFF;

    #10 $display("\n2**912 * 2**111:");
    #10 assign a = 64'h78F0000000000000; assign b = 64'h46E0000000000000;
    #10 assign a = 64'h78FFFFFFFFFFFFFF; assign b = 64'h46EFFFFFFFFFFFFF;

    #10 $display("\n2**913 * 2**110:");
    #10 assign a = 64'h7900000000000000; assign b = 64'h46D0000000000000;
    #10 assign a = 64'h790FFFFFFFFFFFFF; assign b = 64'h46DFFFFFFFFFFFFF;

    #10 $display("\n2**914 * 2**109:");
    #10 assign a = 64'h7910000000000000; assign b = 64'h46C0000000000000;
    #10 assign a = 64'h791FFFFFFFFFFFFF; assign b = 64'h46CFFFFFFFFFFFFF;

    #10 $display("\n2**915 * 2**108:");
    #10 assign a = 64'h7920000000000000; assign b = 64'h46B0000000000000;
    #10 assign a = 64'h792FFFFFFFFFFFFF; assign b = 64'h46BFFFFFFFFFFFFF;

    #10 $display("\n2**916 * 2**107:");
    #10 assign a = 64'h7930000000000000; assign b = 64'h46A0000000000000;
    #10 assign a = 64'h793FFFFFFFFFFFFF; assign b = 64'h46AFFFFFFFFFFFFF;

    #10 $display("\n2**917 * 2**106:");
    #10 assign a = 64'h7940000000000000; assign b = 64'h4690000000000000;
    #10 assign a = 64'h794FFFFFFFFFFFFF; assign b = 64'h469FFFFFFFFFFFFF;

    #10 $display("\n2**918 * 2**105:");
    #10 assign a = 64'h7950000000000000; assign b = 64'h4680000000000000;
    #10 assign a = 64'h795FFFFFFFFFFFFF; assign b = 64'h468FFFFFFFFFFFFF;

    #10 $display("\n2**919 * 2**104:");
    #10 assign a = 64'h7960000000000000; assign b = 64'h4670000000000000;
    #10 assign a = 64'h796FFFFFFFFFFFFF; assign b = 64'h467FFFFFFFFFFFFF;

    #10 $display("\n2**920 * 2**103:");
    #10 assign a = 64'h7970000000000000; assign b = 64'h4660000000000000;
    #10 assign a = 64'h797FFFFFFFFFFFFF; assign b = 64'h466FFFFFFFFFFFFF;

    #10 $display("\n2**921 * 2**102:");
    #10 assign a = 64'h7980000000000000; assign b = 64'h4650000000000000;
    #10 assign a = 64'h798FFFFFFFFFFFFF; assign b = 64'h465FFFFFFFFFFFFF;

    #10 $display("\n2**922 * 2**101:");
    #10 assign a = 64'h7990000000000000; assign b = 64'h4640000000000000;
    #10 assign a = 64'h799FFFFFFFFFFFFF; assign b = 64'h464FFFFFFFFFFFFF;

    #10 $display("\n2**923 * 2**100:");
    #10 assign a = 64'h79A0000000000000; assign b = 64'h4630000000000000;
    #10 assign a = 64'h79AFFFFFFFFFFFFF; assign b = 64'h463FFFFFFFFFFFFF;

    #10 $display("\n2**924 * 2**99:");
    #10 assign a = 64'h79B0000000000000; assign b = 64'h4620000000000000;
    #10 assign a = 64'h79BFFFFFFFFFFFFF; assign b = 64'h462FFFFFFFFFFFFF;

    #10 $display("\n2**925 * 2**98:");
    #10 assign a = 64'h79C0000000000000; assign b = 64'h4610000000000000;
    #10 assign a = 64'h79CFFFFFFFFFFFFF; assign b = 64'h461FFFFFFFFFFFFF;

    #10 $display("\n2**926 * 2**97:");
    #10 assign a = 64'h79D0000000000000; assign b = 64'h4600000000000000;
    #10 assign a = 64'h79DFFFFFFFFFFFFF; assign b = 64'h460FFFFFFFFFFFFF;

    #10 $display("\n2**927 * 2**96:");
    #10 assign a = 64'h79E0000000000000; assign b = 64'h45F0000000000000;
    #10 assign a = 64'h79EFFFFFFFFFFFFF; assign b = 64'h45FFFFFFFFFFFFFF;

    #10 $display("\n2**928 * 2**95:");
    #10 assign a = 64'h79F0000000000000; assign b = 64'h45E0000000000000;
    #10 assign a = 64'h79FFFFFFFFFFFFFF; assign b = 64'h45EFFFFFFFFFFFFF;

    #10 $display("\n2**929 * 2**94:");
    #10 assign a = 64'h7A00000000000000; assign b = 64'h45D0000000000000;
    #10 assign a = 64'h7A0FFFFFFFFFFFFF; assign b = 64'h45DFFFFFFFFFFFFF;

    #10 $display("\n2**930 * 2**93:");
    #10 assign a = 64'h7A10000000000000; assign b = 64'h45C0000000000000;
    #10 assign a = 64'h7A1FFFFFFFFFFFFF; assign b = 64'h45CFFFFFFFFFFFFF;

    #10 $display("\n2**931 * 2**92:");
    #10 assign a = 64'h7A20000000000000; assign b = 64'h45B0000000000000;
    #10 assign a = 64'h7A2FFFFFFFFFFFFF; assign b = 64'h45BFFFFFFFFFFFFF;

    #10 $display("\n2**932 * 2**91:");
    #10 assign a = 64'h7A30000000000000; assign b = 64'h45A0000000000000;
    #10 assign a = 64'h7A3FFFFFFFFFFFFF; assign b = 64'h45AFFFFFFFFFFFFF;

    #10 $display("\n2**933 * 2**90:");
    #10 assign a = 64'h7A40000000000000; assign b = 64'h4590000000000000;
    #10 assign a = 64'h7A4FFFFFFFFFFFFF; assign b = 64'h459FFFFFFFFFFFFF;

    #10 $display("\n2**934 * 2**89:");
    #10 assign a = 64'h7A50000000000000; assign b = 64'h4580000000000000;
    #10 assign a = 64'h7A5FFFFFFFFFFFFF; assign b = 64'h458FFFFFFFFFFFFF;

    #10 $display("\n2**935 * 2**88:");
    #10 assign a = 64'h7A60000000000000; assign b = 64'h4570000000000000;
    #10 assign a = 64'h7A6FFFFFFFFFFFFF; assign b = 64'h457FFFFFFFFFFFFF;

    #10 $display("\n2**936 * 2**87:");
    #10 assign a = 64'h7A70000000000000; assign b = 64'h4560000000000000;
    #10 assign a = 64'h7A7FFFFFFFFFFFFF; assign b = 64'h456FFFFFFFFFFFFF;

    #10 $display("\n2**937 * 2**86:");
    #10 assign a = 64'h7A80000000000000; assign b = 64'h4550000000000000;
    #10 assign a = 64'h7A8FFFFFFFFFFFFF; assign b = 64'h455FFFFFFFFFFFFF;

    #10 $display("\n2**938 * 2**85:");
    #10 assign a = 64'h7A90000000000000; assign b = 64'h4540000000000000;
    #10 assign a = 64'h7A9FFFFFFFFFFFFF; assign b = 64'h454FFFFFFFFFFFFF;

    #10 $display("\n2**939 * 2**84:");
    #10 assign a = 64'h7AA0000000000000; assign b = 64'h4530000000000000;
    #10 assign a = 64'h7AAFFFFFFFFFFFFF; assign b = 64'h453FFFFFFFFFFFFF;

    #10 $display("\n2**940 * 2**83:");
    #10 assign a = 64'h7AB0000000000000; assign b = 64'h4520000000000000;
    #10 assign a = 64'h7ABFFFFFFFFFFFFF; assign b = 64'h452FFFFFFFFFFFFF;

    #10 $display("\n2**941 * 2**82:");
    #10 assign a = 64'h7AC0000000000000; assign b = 64'h4510000000000000;
    #10 assign a = 64'h7ACFFFFFFFFFFFFF; assign b = 64'h451FFFFFFFFFFFFF;

    #10 $display("\n2**942 * 2**81:");
    #10 assign a = 64'h7AD0000000000000; assign b = 64'h4500000000000000;
    #10 assign a = 64'h7ADFFFFFFFFFFFFF; assign b = 64'h450FFFFFFFFFFFFF;

    #10 $display("\n2**943 * 2**80:");
    #10 assign a = 64'h7AE0000000000000; assign b = 64'h44F0000000000000;
    #10 assign a = 64'h7AEFFFFFFFFFFFFF; assign b = 64'h44FFFFFFFFFFFFFF;

    #10 $display("\n2**944 * 2**79:");
    #10 assign a = 64'h7AF0000000000000; assign b = 64'h44E0000000000000;
    #10 assign a = 64'h7AFFFFFFFFFFFFFF; assign b = 64'h44EFFFFFFFFFFFFF;

    #10 $display("\n2**945 * 2**78:");
    #10 assign a = 64'h7B00000000000000; assign b = 64'h44D0000000000000;
    #10 assign a = 64'h7B0FFFFFFFFFFFFF; assign b = 64'h44DFFFFFFFFFFFFF;

    #10 $display("\n2**946 * 2**77:");
    #10 assign a = 64'h7B10000000000000; assign b = 64'h44C0000000000000;
    #10 assign a = 64'h7B1FFFFFFFFFFFFF; assign b = 64'h44CFFFFFFFFFFFFF;

    #10 $display("\n2**947 * 2**76:");
    #10 assign a = 64'h7B20000000000000; assign b = 64'h44B0000000000000;
    #10 assign a = 64'h7B2FFFFFFFFFFFFF; assign b = 64'h44BFFFFFFFFFFFFF;

    #10 $display("\n2**948 * 2**75:");
    #10 assign a = 64'h7B30000000000000; assign b = 64'h44A0000000000000;
    #10 assign a = 64'h7B3FFFFFFFFFFFFF; assign b = 64'h44AFFFFFFFFFFFFF;

    #10 $display("\n2**949 * 2**74:");
    #10 assign a = 64'h7B40000000000000; assign b = 64'h4490000000000000;
    #10 assign a = 64'h7B4FFFFFFFFFFFFF; assign b = 64'h449FFFFFFFFFFFFF;

    #10 $display("\n2**950 * 2**73:");
    #10 assign a = 64'h7B50000000000000; assign b = 64'h4480000000000000;
    #10 assign a = 64'h7B5FFFFFFFFFFFFF; assign b = 64'h448FFFFFFFFFFFFF;

    #10 $display("\n2**951 * 2**72:");
    #10 assign a = 64'h7B60000000000000; assign b = 64'h4470000000000000;
    #10 assign a = 64'h7B6FFFFFFFFFFFFF; assign b = 64'h447FFFFFFFFFFFFF;

    #10 $display("\n2**952 * 2**71:");
    #10 assign a = 64'h7B70000000000000; assign b = 64'h4460000000000000;
    #10 assign a = 64'h7B7FFFFFFFFFFFFF; assign b = 64'h446FFFFFFFFFFFFF;

    #10 $display("\n2**953 * 2**70:");
    #10 assign a = 64'h7B80000000000000; assign b = 64'h4450000000000000;
    #10 assign a = 64'h7B8FFFFFFFFFFFFF; assign b = 64'h445FFFFFFFFFFFFF;

    #10 $display("\n2**954 * 2**69:");
    #10 assign a = 64'h7B90000000000000; assign b = 64'h4440000000000000;
    #10 assign a = 64'h7B9FFFFFFFFFFFFF; assign b = 64'h444FFFFFFFFFFFFF;

    #10 $display("\n2**955 * 2**68:");
    #10 assign a = 64'h7BA0000000000000; assign b = 64'h4430000000000000;
    #10 assign a = 64'h7BAFFFFFFFFFFFFF; assign b = 64'h443FFFFFFFFFFFFF;

    #10 $display("\n2**956 * 2**67:");
    #10 assign a = 64'h7BB0000000000000; assign b = 64'h4420000000000000;
    #10 assign a = 64'h7BBFFFFFFFFFFFFF; assign b = 64'h442FFFFFFFFFFFFF;

    #10 $display("\n2**957 * 2**66:");
    #10 assign a = 64'h7BC0000000000000; assign b = 64'h4410000000000000;
    #10 assign a = 64'h7BCFFFFFFFFFFFFF; assign b = 64'h441FFFFFFFFFFFFF;

    #10 $display("\n2**958 * 2**65:");
    #10 assign a = 64'h7BD0000000000000; assign b = 64'h4400000000000000;
    #10 assign a = 64'h7BDFFFFFFFFFFFFF; assign b = 64'h440FFFFFFFFFFFFF;

    #10 $display("\n2**959 * 2**64:");
    #10 assign a = 64'h7BE0000000000000; assign b = 64'h43F0000000000000;
    #10 assign a = 64'h7BEFFFFFFFFFFFFF; assign b = 64'h43FFFFFFFFFFFFFF;

    #10 $display("\n2**960 * 2**63:");
    #10 assign a = 64'h7BF0000000000000; assign b = 64'h43E0000000000000;
    #10 assign a = 64'h7BFFFFFFFFFFFFFF; assign b = 64'h43EFFFFFFFFFFFFF;

    #10 $display("\n2**961 * 2**62:");
    #10 assign a = 64'h7C00000000000000; assign b = 64'h43D0000000000000;
    #10 assign a = 64'h7C0FFFFFFFFFFFFF; assign b = 64'h43DFFFFFFFFFFFFF;

    #10 $display("\n2**962 * 2**61:");
    #10 assign a = 64'h7C10000000000000; assign b = 64'h43C0000000000000;
    #10 assign a = 64'h7C1FFFFFFFFFFFFF; assign b = 64'h43CFFFFFFFFFFFFF;

    #10 $display("\n2**963 * 2**60:");
    #10 assign a = 64'h7C20000000000000; assign b = 64'h43B0000000000000;
    #10 assign a = 64'h7C2FFFFFFFFFFFFF; assign b = 64'h43BFFFFFFFFFFFFF;

    #10 $display("\n2**964 * 2**59:");
    #10 assign a = 64'h7C30000000000000; assign b = 64'h43A0000000000000;
    #10 assign a = 64'h7C3FFFFFFFFFFFFF; assign b = 64'h43AFFFFFFFFFFFFF;

    #10 $display("\n2**965 * 2**58:");
    #10 assign a = 64'h7C40000000000000; assign b = 64'h4390000000000000;
    #10 assign a = 64'h7C4FFFFFFFFFFFFF; assign b = 64'h439FFFFFFFFFFFFF;

    #10 $display("\n2**966 * 2**57:");
    #10 assign a = 64'h7C50000000000000; assign b = 64'h4380000000000000;
    #10 assign a = 64'h7C5FFFFFFFFFFFFF; assign b = 64'h438FFFFFFFFFFFFF;

    #10 $display("\n2**967 * 2**56:");
    #10 assign a = 64'h7C60000000000000; assign b = 64'h4370000000000000;
    #10 assign a = 64'h7C6FFFFFFFFFFFFF; assign b = 64'h437FFFFFFFFFFFFF;

    #10 $display("\n2**968 * 2**55:");
    #10 assign a = 64'h7C70000000000000; assign b = 64'h4360000000000000;
    #10 assign a = 64'h7C7FFFFFFFFFFFFF; assign b = 64'h436FFFFFFFFFFFFF;

    #10 $display("\n2**969 * 2**54:");
    #10 assign a = 64'h7C80000000000000; assign b = 64'h4350000000000000;
    #10 assign a = 64'h7C8FFFFFFFFFFFFF; assign b = 64'h435FFFFFFFFFFFFF;

    #10 $display("\n2**970 * 2**53:");
    #10 assign a = 64'h7C90000000000000; assign b = 64'h4340000000000000;
    #10 assign a = 64'h7C9FFFFFFFFFFFFF; assign b = 64'h434FFFFFFFFFFFFF;

    #10 $display("\n2**971 * 2**52:");
    #10 assign a = 64'h7CA0000000000000; assign b = 64'h4330000000000000;
    #10 assign a = 64'h7CAFFFFFFFFFFFFF; assign b = 64'h433FFFFFFFFFFFFF;

    #10 $display("\n2**972 * 2**51:");
    #10 assign a = 64'h7CB0000000000000; assign b = 64'h4320000000000000;
    #10 assign a = 64'h7CBFFFFFFFFFFFFF; assign b = 64'h432FFFFFFFFFFFFF;

    #10 $display("\n2**973 * 2**50:");
    #10 assign a = 64'h7CC0000000000000; assign b = 64'h4310000000000000;
    #10 assign a = 64'h7CCFFFFFFFFFFFFF; assign b = 64'h431FFFFFFFFFFFFF;

    #10 $display("\n2**974 * 2**49:");
    #10 assign a = 64'h7CD0000000000000; assign b = 64'h4300000000000000;
    #10 assign a = 64'h7CDFFFFFFFFFFFFF; assign b = 64'h430FFFFFFFFFFFFF;

    #10 $display("\n2**975 * 2**48:");
    #10 assign a = 64'h7CE0000000000000; assign b = 64'h42F0000000000000;
    #10 assign a = 64'h7CEFFFFFFFFFFFFF; assign b = 64'h42FFFFFFFFFFFFFF;

    #10 $display("\n2**976 * 2**47:");
    #10 assign a = 64'h7CF0000000000000; assign b = 64'h42E0000000000000;
    #10 assign a = 64'h7CFFFFFFFFFFFFFF; assign b = 64'h42EFFFFFFFFFFFFF;

    #10 $display("\n2**977 * 2**46:");
    #10 assign a = 64'h7D00000000000000; assign b = 64'h42D0000000000000;
    #10 assign a = 64'h7D0FFFFFFFFFFFFF; assign b = 64'h42DFFFFFFFFFFFFF;

    #10 $display("\n2**978 * 2**45:");
    #10 assign a = 64'h7D10000000000000; assign b = 64'h42C0000000000000;
    #10 assign a = 64'h7D1FFFFFFFFFFFFF; assign b = 64'h42CFFFFFFFFFFFFF;

    #10 $display("\n2**979 * 2**44:");
    #10 assign a = 64'h7D20000000000000; assign b = 64'h42B0000000000000;
    #10 assign a = 64'h7D2FFFFFFFFFFFFF; assign b = 64'h42BFFFFFFFFFFFFF;

    #10 $display("\n2**980 * 2**43:");
    #10 assign a = 64'h7D30000000000000; assign b = 64'h42A0000000000000;
    #10 assign a = 64'h7D3FFFFFFFFFFFFF; assign b = 64'h42AFFFFFFFFFFFFF;

    #10 $display("\n2**981 * 2**42:");
    #10 assign a = 64'h7D40000000000000; assign b = 64'h4290000000000000;
    #10 assign a = 64'h7D4FFFFFFFFFFFFF; assign b = 64'h429FFFFFFFFFFFFF;

    #10 $display("\n2**982 * 2**41:");
    #10 assign a = 64'h7D50000000000000; assign b = 64'h4280000000000000;
    #10 assign a = 64'h7D5FFFFFFFFFFFFF; assign b = 64'h428FFFFFFFFFFFFF;

    #10 $display("\n2**983 * 2**40:");
    #10 assign a = 64'h7D60000000000000; assign b = 64'h4270000000000000;
    #10 assign a = 64'h7D6FFFFFFFFFFFFF; assign b = 64'h427FFFFFFFFFFFFF;

    #10 $display("\n2**984 * 2**39:");
    #10 assign a = 64'h7D70000000000000; assign b = 64'h4260000000000000;
    #10 assign a = 64'h7D7FFFFFFFFFFFFF; assign b = 64'h426FFFFFFFFFFFFF;

    #10 $display("\n2**985 * 2**38:");
    #10 assign a = 64'h7D80000000000000; assign b = 64'h4250000000000000;
    #10 assign a = 64'h7D8FFFFFFFFFFFFF; assign b = 64'h425FFFFFFFFFFFFF;

    #10 $display("\n2**986 * 2**37:");
    #10 assign a = 64'h7D90000000000000; assign b = 64'h4240000000000000;
    #10 assign a = 64'h7D9FFFFFFFFFFFFF; assign b = 64'h424FFFFFFFFFFFFF;

    #10 $display("\n2**987 * 2**36:");
    #10 assign a = 64'h7DA0000000000000; assign b = 64'h4230000000000000;
    #10 assign a = 64'h7DAFFFFFFFFFFFFF; assign b = 64'h423FFFFFFFFFFFFF;

    #10 $display("\n2**988 * 2**35:");
    #10 assign a = 64'h7DB0000000000000; assign b = 64'h4220000000000000;
    #10 assign a = 64'h7DBFFFFFFFFFFFFF; assign b = 64'h422FFFFFFFFFFFFF;

    #10 $display("\n2**989 * 2**34:");
    #10 assign a = 64'h7DC0000000000000; assign b = 64'h4210000000000000;
    #10 assign a = 64'h7DCFFFFFFFFFFFFF; assign b = 64'h421FFFFFFFFFFFFF;

    #10 $display("\n2**990 * 2**33:");
    #10 assign a = 64'h7DD0000000000000; assign b = 64'h4200000000000000;
    #10 assign a = 64'h7DDFFFFFFFFFFFFF; assign b = 64'h420FFFFFFFFFFFFF;

    #10 $display("\n2**991 * 2**32:");
    #10 assign a = 64'h7DE0000000000000; assign b = 64'h41F0000000000000;
    #10 assign a = 64'h7DEFFFFFFFFFFFFF; assign b = 64'h41FFFFFFFFFFFFFF;

    #10 $display("\n2**992 * 2**31:");
    #10 assign a = 64'h7DF0000000000000; assign b = 64'h41E0000000000000;
    #10 assign a = 64'h7DFFFFFFFFFFFFFF; assign b = 64'h41EFFFFFFFFFFFFF;

    #10 $display("\n2**993 * 2**30:");
    #10 assign a = 64'h7E00000000000000; assign b = 64'h41D0000000000000;
    #10 assign a = 64'h7E0FFFFFFFFFFFFF; assign b = 64'h41DFFFFFFFFFFFFF;

    #10 $display("\n2**994 * 2**29:");
    #10 assign a = 64'h7E10000000000000; assign b = 64'h41C0000000000000;
    #10 assign a = 64'h7E1FFFFFFFFFFFFF; assign b = 64'h41CFFFFFFFFFFFFF;

    #10 $display("\n2**995 * 2**28:");
    #10 assign a = 64'h7E20000000000000; assign b = 64'h41B0000000000000;
    #10 assign a = 64'h7E2FFFFFFFFFFFFF; assign b = 64'h41BFFFFFFFFFFFFF;

    #10 $display("\n2**996 * 2**27:");
    #10 assign a = 64'h7E30000000000000; assign b = 64'h41A0000000000000;
    #10 assign a = 64'h7E3FFFFFFFFFFFFF; assign b = 64'h41AFFFFFFFFFFFFF;

    #10 $display("\n2**997 * 2**26:");
    #10 assign a = 64'h7E40000000000000; assign b = 64'h4190000000000000;
    #10 assign a = 64'h7E4FFFFFFFFFFFFF; assign b = 64'h419FFFFFFFFFFFFF;

    #10 $display("\n2**998 * 2**25:");
    #10 assign a = 64'h7E50000000000000; assign b = 64'h4180000000000000;
    #10 assign a = 64'h7E5FFFFFFFFFFFFF; assign b = 64'h418FFFFFFFFFFFFF;

    #10 $display("\n2**999 * 2**24:");
    #10 assign a = 64'h7E60000000000000; assign b = 64'h4170000000000000;
    #10 assign a = 64'h7E6FFFFFFFFFFFFF; assign b = 64'h417FFFFFFFFFFFFF;

    #10 $display("\n2**1000 * 2**23:");
    #10 assign a = 64'h7E70000000000000; assign b = 64'h4160000000000000;
    #10 assign a = 64'h7E7FFFFFFFFFFFFF; assign b = 64'h416FFFFFFFFFFFFF;

    #10 $display("\n2**1001 * 2**22:");
    #10 assign a = 64'h7E80000000000000; assign b = 64'h4150000000000000;
    #10 assign a = 64'h7E8FFFFFFFFFFFFF; assign b = 64'h415FFFFFFFFFFFFF;

    #10 $display("\n2**1002 * 2**21:");
    #10 assign a = 64'h7E90000000000000; assign b = 64'h4140000000000000;
    #10 assign a = 64'h7E9FFFFFFFFFFFFF; assign b = 64'h414FFFFFFFFFFFFF;

    #10 $display("\n2**1003 * 2**20:");
    #10 assign a = 64'h7EA0000000000000; assign b = 64'h4130000000000000;
    #10 assign a = 64'h7EAFFFFFFFFFFFFF; assign b = 64'h413FFFFFFFFFFFFF;

    #10 $display("\n2**1004 * 2**19:");
    #10 assign a = 64'h7EB0000000000000; assign b = 64'h4120000000000000;
    #10 assign a = 64'h7EBFFFFFFFFFFFFF; assign b = 64'h412FFFFFFFFFFFFF;

    #10 $display("\n2**1005 * 2**18:");
    #10 assign a = 64'h7EC0000000000000; assign b = 64'h4110000000000000;
    #10 assign a = 64'h7ECFFFFFFFFFFFFF; assign b = 64'h411FFFFFFFFFFFFF;

    #10 $display("\n2**1006 * 2**17:");
    #10 assign a = 64'h7ED0000000000000; assign b = 64'h4100000000000000;
    #10 assign a = 64'h7EDFFFFFFFFFFFFF; assign b = 64'h410FFFFFFFFFFFFF;

    #10 $display("\n2**1007 * 2**16:");
    #10 assign a = 64'h7EE0000000000000; assign b = 64'h40F0000000000000;
    #10 assign a = 64'h7EEFFFFFFFFFFFFF; assign b = 64'h40FFFFFFFFFFFFFF;

    #10 $display("\n2**1008 * 2**15:");
    #10 assign a = 64'h7EF0000000000000; assign b = 64'h40E0000000000000;
    #10 assign a = 64'h7EFFFFFFFFFFFFFF; assign b = 64'h40EFFFFFFFFFFFFF;

    #10 $display("\n2**1009 * 2**14:");
    #10 assign a = 64'h7F00000000000000; assign b = 64'h40D0000000000000;
    #10 assign a = 64'h7F0FFFFFFFFFFFFF; assign b = 64'h40DFFFFFFFFFFFFF;

    #10 $display("\n2**1010 * 2**13:");
    #10 assign a = 64'h7F10000000000000; assign b = 64'h40C0000000000000;
    #10 assign a = 64'h7F1FFFFFFFFFFFFF; assign b = 64'h40CFFFFFFFFFFFFF;

    #10 $display("\n2**1011 * 2**12:");
    #10 assign a = 64'h7F20000000000000; assign b = 64'h40B0000000000000;
    #10 assign a = 64'h7F2FFFFFFFFFFFFF; assign b = 64'h40BFFFFFFFFFFFFF;

    #10 $display("\n2**1012 * 2**11:");
    #10 assign a = 64'h7F30000000000000; assign b = 64'h40A0000000000000;
    #10 assign a = 64'h7F3FFFFFFFFFFFFF; assign b = 64'h40AFFFFFFFFFFFFF;

    #10 $display("\n2**1013 * 2**10:");
    #10 assign a = 64'h7F40000000000000; assign b = 64'h4090000000000000;
    #10 assign a = 64'h7F4FFFFFFFFFFFFF; assign b = 64'h409FFFFFFFFFFFFF;

    #10 $display("\n2**1014 * 2**9:");
    #10 assign a = 64'h7F50000000000000; assign b = 64'h4080000000000000;
    #10 assign a = 64'h7F5FFFFFFFFFFFFF; assign b = 64'h408FFFFFFFFFFFFF;

    #10 $display("\n2**1015 * 2**8:");
    #10 assign a = 64'h7F60000000000000; assign b = 64'h4070000000000000;
    #10 assign a = 64'h7F6FFFFFFFFFFFFF; assign b = 64'h407FFFFFFFFFFFFF;

    #10 $display("\n2**1016 * 2**7:");
    #10 assign a = 64'h7F70000000000000; assign b = 64'h4060000000000000;
    #10 assign a = 64'h7F7FFFFFFFFFFFFF; assign b = 64'h406FFFFFFFFFFFFF;

    #10 $display("\n2**1017 * 2**6:");
    #10 assign a = 64'h7F80000000000000; assign b = 64'h4050000000000000;
    #10 assign a = 64'h7F8FFFFFFFFFFFFF; assign b = 64'h405FFFFFFFFFFFFF;

    #10 $display("\n2**1018 * 2**5:");
    #10 assign a = 64'h7F90000000000000; assign b = 64'h4040000000000000;
    #10 assign a = 64'h7F9FFFFFFFFFFFFF; assign b = 64'h404FFFFFFFFFFFFF;

    #10 $display("\n2**1019 * 2**4:");
    #10 assign a = 64'h7FA0000000000000; assign b = 64'h4030000000000000;
    #10 assign a = 64'h7FAFFFFFFFFFFFFF; assign b = 64'h403FFFFFFFFFFFFF;

    #10 $display("\n2**1020 * 2**3:");
    #10 assign a = 64'h7FB0000000000000; assign b = 64'h4020000000000000;
    #10 assign a = 64'h7FBFFFFFFFFFFFFF; assign b = 64'h402FFFFFFFFFFFFF;

    #10 $display("\n2**1021 * 2**2:");
    #10 assign a = 64'h7FC0000000000000; assign b = 64'h4010000000000000;
    #10 assign a = 64'h7FCFFFFFFFFFFFFF; assign b = 64'h401FFFFFFFFFFFFF;

    #10 $display("\n2**1022 * 2**1:");
    #10 assign a = 64'h7FD0000000000000; assign b = 64'h4000000000000000;
    #10 assign a = 64'h7FDFFFFFFFFFFFFF; assign b = 64'h400FFFFFFFFFFFFF;

    #10 $display("\n2**1023 * 2**0:");
    #10 assign a = 64'h7FE0000000000000; assign b = 64'h3FF0000000000000;
    #10 assign a = 64'h7FEFFFFFFFFFFFFF; assign b = 64'h3FFFFFFFFFFFFFFF;

    #10 $display("\n2**-1074 * 2**51:");
    #10 assign a = 64'h0000000000000001; assign b = 64'h4320000000000000;
    #10 assign a = 64'h0000000000000001; assign b = 64'h432FFFFFFFFFFFFF;

    #10 $display("\n2**-1073 * 2**50:");
    #10 assign a = 64'h0000000000000002; assign b = 64'h4310000000000000;
    #10 assign a = 64'h0000000000000003; assign b = 64'h431FFFFFFFFFFFFF;

    #10 $display("\n2**-1072 * 2**49:");
    #10 assign a = 64'h0000000000000004; assign b = 64'h4300000000000000;
    #10 assign a = 64'h0000000000000007; assign b = 64'h430FFFFFFFFFFFFF;

    #10 $display("\n2**-1071 * 2**48:");
    #10 assign a = 64'h0000000000000008; assign b = 64'h42F0000000000000;
    #10 assign a = 64'h000000000000000F; assign b = 64'h42FFFFFFFFFFFFFF;

    #10 $display("\n2**-1070 * 2**47:");
    #10 assign a = 64'h0000000000000010; assign b = 64'h42E0000000000000;
    #10 assign a = 64'h000000000000001F; assign b = 64'h42EFFFFFFFFFFFFF;

    #10 $display("\n2**-1069 * 2**46:");
    #10 assign a = 64'h0000000000000020; assign b = 64'h42D0000000000000;
    #10 assign a = 64'h000000000000003F; assign b = 64'h42DFFFFFFFFFFFFF;

    #10 $display("\n2**-1068 * 2**45:");
    #10 assign a = 64'h0000000000000040; assign b = 64'h42C0000000000000;
    #10 assign a = 64'h000000000000007F; assign b = 64'h42CFFFFFFFFFFFFF;

    #10 $display("\n2**-1067 * 2**44:");
    #10 assign a = 64'h0000000000000080; assign b = 64'h42B0000000000000;
    #10 assign a = 64'h00000000000000FF; assign b = 64'h42BFFFFFFFFFFFFF;

    #10 $display("\n2**-1066 * 2**43:");
    #10 assign a = 64'h0000000000000100; assign b = 64'h42A0000000000000;
    #10 assign a = 64'h00000000000001FF; assign b = 64'h42AFFFFFFFFFFFFF;

    #10 $display("\n2**-1065 * 2**42:");
    #10 assign a = 64'h0000000000000200; assign b = 64'h4290000000000000;
    #10 assign a = 64'h00000000000003FF; assign b = 64'h429FFFFFFFFFFFFF;

    #10 $display("\n2**-1064 * 2**41:");
    #10 assign a = 64'h0000000000000400; assign b = 64'h4280000000000000;
    #10 assign a = 64'h00000000000007FF; assign b = 64'h428FFFFFFFFFFFFF;

    #10 $display("\n2**-1063 * 2**40:");
    #10 assign a = 64'h0000000000000800; assign b = 64'h4270000000000000;
    #10 assign a = 64'h0000000000000FFF; assign b = 64'h427FFFFFFFFFFFFF;

    #10 $display("\n2**-1062 * 2**39:");
    #10 assign a = 64'h0000000000001000; assign b = 64'h4260000000000000;
    #10 assign a = 64'h0000000000001FFF; assign b = 64'h426FFFFFFFFFFFFF;

    #10 $display("\n2**-1061 * 2**38:");
    #10 assign a = 64'h0000000000002000; assign b = 64'h4250000000000000;
    #10 assign a = 64'h0000000000003FFF; assign b = 64'h425FFFFFFFFFFFFF;

    #10 $display("\n2**-1060 * 2**37:");
    #10 assign a = 64'h0000000000004000; assign b = 64'h4240000000000000;
    #10 assign a = 64'h0000000000007FFF; assign b = 64'h424FFFFFFFFFFFFF;

    #10 $display("\n2**-1059 * 2**36:");
    #10 assign a = 64'h0000000000008000; assign b = 64'h4230000000000000;
    #10 assign a = 64'h000000000000FFFF; assign b = 64'h423FFFFFFFFFFFFF;

    #10 $display("\n2**-1058 * 2**35:");
    #10 assign a = 64'h0000000000010000; assign b = 64'h4220000000000000;
    #10 assign a = 64'h000000000001FFFF; assign b = 64'h422FFFFFFFFFFFFF;

    #10 $display("\n2**-1057 * 2**34:");
    #10 assign a = 64'h0000000000020000; assign b = 64'h4210000000000000;
    #10 assign a = 64'h000000000003FFFF; assign b = 64'h421FFFFFFFFFFFFF;

    #10 $display("\n2**-1056 * 2**33:");
    #10 assign a = 64'h0000000000040000; assign b = 64'h4200000000000000;
    #10 assign a = 64'h000000000007FFFF; assign b = 64'h420FFFFFFFFFFFFF;

    #10 $display("\n2**-1055 * 2**32:");
    #10 assign a = 64'h0000000000080000; assign b = 64'h41F0000000000000;
    #10 assign a = 64'h00000000000FFFFF; assign b = 64'h41FFFFFFFFFFFFFF;

    #10 $display("\n2**-1054 * 2**31:");
    #10 assign a = 64'h0000000000100000; assign b = 64'h41E0000000000000;
    #10 assign a = 64'h00000000001FFFFF; assign b = 64'h41EFFFFFFFFFFFFF;

    #10 $display("\n2**-1053 * 2**30:");
    #10 assign a = 64'h0000000000200000; assign b = 64'h41D0000000000000;
    #10 assign a = 64'h00000000003FFFFF; assign b = 64'h41DFFFFFFFFFFFFF;

    #10 $display("\n2**-1052 * 2**29:");
    #10 assign a = 64'h0000000000400000; assign b = 64'h41C0000000000000;
    #10 assign a = 64'h00000000007FFFFF; assign b = 64'h41CFFFFFFFFFFFFF;

    #10 $display("\n2**-1051 * 2**28:");
    #10 assign a = 64'h0000000000800000; assign b = 64'h41B0000000000000;
    #10 assign a = 64'h0000000000FFFFFF; assign b = 64'h41BFFFFFFFFFFFFF;

    #10 $display("\n2**-1050 * 2**27:");
    #10 assign a = 64'h0000000001000000; assign b = 64'h41A0000000000000;
    #10 assign a = 64'h0000000001FFFFFF; assign b = 64'h41AFFFFFFFFFFFFF;

    #10 $display("\n2**-1049 * 2**26:");
    #10 assign a = 64'h0000000002000000; assign b = 64'h4190000000000000;
    #10 assign a = 64'h0000000003FFFFFF; assign b = 64'h419FFFFFFFFFFFFF;

    #10 $display("\n2**-1048 * 2**25:");
    #10 assign a = 64'h0000000004000000; assign b = 64'h4180000000000000;
    #10 assign a = 64'h0000000007FFFFFF; assign b = 64'h418FFFFFFFFFFFFF;

    #10 $display("\n2**-1047 * 2**24:");
    #10 assign a = 64'h0000000008000000; assign b = 64'h4170000000000000;
    #10 assign a = 64'h000000000FFFFFFF; assign b = 64'h417FFFFFFFFFFFFF;

    #10 $display("\n2**-1046 * 2**23:");
    #10 assign a = 64'h0000000010000000; assign b = 64'h4160000000000000;
    #10 assign a = 64'h000000001FFFFFFF; assign b = 64'h416FFFFFFFFFFFFF;

    #10 $display("\n2**-1045 * 2**22:");
    #10 assign a = 64'h0000000020000000; assign b = 64'h4150000000000000;
    #10 assign a = 64'h000000003FFFFFFF; assign b = 64'h415FFFFFFFFFFFFF;

    #10 $display("\n2**-1044 * 2**21:");
    #10 assign a = 64'h0000000040000000; assign b = 64'h4140000000000000;
    #10 assign a = 64'h000000007FFFFFFF; assign b = 64'h414FFFFFFFFFFFFF;

    #10 $display("\n2**-1043 * 2**20:");
    #10 assign a = 64'h0000000080000000; assign b = 64'h4130000000000000;
    #10 assign a = 64'h00000000FFFFFFFF; assign b = 64'h413FFFFFFFFFFFFF;

    #10 $display("\n2**-1042 * 2**19:");
    #10 assign a = 64'h0000000100000000; assign b = 64'h4120000000000000;
    #10 assign a = 64'h00000001FFFFFFFF; assign b = 64'h412FFFFFFFFFFFFF;

    #10 $display("\n2**-1041 * 2**18:");
    #10 assign a = 64'h0000000200000000; assign b = 64'h4110000000000000;
    #10 assign a = 64'h00000003FFFFFFFF; assign b = 64'h411FFFFFFFFFFFFF;

    #10 $display("\n2**-1040 * 2**17:");
    #10 assign a = 64'h0000000400000000; assign b = 64'h4100000000000000;
    #10 assign a = 64'h00000007FFFFFFFF; assign b = 64'h410FFFFFFFFFFFFF;

    #10 $display("\n2**-1039 * 2**16:");
    #10 assign a = 64'h0000000800000000; assign b = 64'h40F0000000000000;
    #10 assign a = 64'h0000000FFFFFFFFF; assign b = 64'h40FFFFFFFFFFFFFF;

    #10 $display("\n2**-1038 * 2**15:");
    #10 assign a = 64'h0000001000000000; assign b = 64'h40E0000000000000;
    #10 assign a = 64'h0000001FFFFFFFFF; assign b = 64'h40EFFFFFFFFFFFFF;

    #10 $display("\n2**-1037 * 2**14:");
    #10 assign a = 64'h0000002000000000; assign b = 64'h40D0000000000000;
    #10 assign a = 64'h0000003FFFFFFFFF; assign b = 64'h40DFFFFFFFFFFFFF;

    #10 $display("\n2**-1036 * 2**13:");
    #10 assign a = 64'h0000004000000000; assign b = 64'h40C0000000000000;
    #10 assign a = 64'h0000007FFFFFFFFF; assign b = 64'h40CFFFFFFFFFFFFF;

    #10 $display("\n2**-1035 * 2**12:");
    #10 assign a = 64'h0000008000000000; assign b = 64'h40B0000000000000;
    #10 assign a = 64'h000000FFFFFFFFFF; assign b = 64'h40BFFFFFFFFFFFFF;

    #10 $display("\n2**-1034 * 2**11:");
    #10 assign a = 64'h0000010000000000; assign b = 64'h40A0000000000000;
    #10 assign a = 64'h000001FFFFFFFFFF; assign b = 64'h40AFFFFFFFFFFFFF;

    #10 $display("\n2**-1033 * 2**10:");
    #10 assign a = 64'h0000020000000000; assign b = 64'h4090000000000000;
    #10 assign a = 64'h000003FFFFFFFFFF; assign b = 64'h409FFFFFFFFFFFFF;

    #10 $display("\n2**-1032 * 2**9:");
    #10 assign a = 64'h0000040000000000; assign b = 64'h4080000000000000;
    #10 assign a = 64'h000007FFFFFFFFFF; assign b = 64'h408FFFFFFFFFFFFF;

    #10 $display("\n2**-1031 * 2**8:");
    #10 assign a = 64'h0000080000000000; assign b = 64'h4070000000000000;
    #10 assign a = 64'h00000FFFFFFFFFFF; assign b = 64'h407FFFFFFFFFFFFF;

    #10 $display("\n2**-1030 * 2**7:");
    #10 assign a = 64'h0000100000000000; assign b = 64'h4060000000000000;
    #10 assign a = 64'h00001FFFFFFFFFFF; assign b = 64'h406FFFFFFFFFFFFF;

    #10 $display("\n2**-1029 * 2**6:");
    #10 assign a = 64'h0000200000000000; assign b = 64'h4050000000000000;
    #10 assign a = 64'h00003FFFFFFFFFFF; assign b = 64'h405FFFFFFFFFFFFF;

    #10 $display("\n2**-1028 * 2**5:");
    #10 assign a = 64'h0000400000000000; assign b = 64'h4040000000000000;
    #10 assign a = 64'h00007FFFFFFFFFFF; assign b = 64'h404FFFFFFFFFFFFF;

    #10 $display("\n2**-1027 * 2**4:");
    #10 assign a = 64'h0000800000000000; assign b = 64'h4030000000000000;
    #10 assign a = 64'h0000FFFFFFFFFFFF; assign b = 64'h403FFFFFFFFFFFFF;

    #10 $display("\n2**-1026 * 2**3:");
    #10 assign a = 64'h0001000000000000; assign b = 64'h4020000000000000;
    #10 assign a = 64'h0001FFFFFFFFFFFF; assign b = 64'h402FFFFFFFFFFFFF;

    #10 $display("\n2**-1025 * 2**2:");
    #10 assign a = 64'h0002000000000000; assign b = 64'h4010000000000000;
    #10 assign a = 64'h0003FFFFFFFFFFFF; assign b = 64'h401FFFFFFFFFFFFF;

    #10 $display("\n2**-1024 * 2**1:");
    #10 assign a = 64'h0004000000000000; assign b = 64'h4000000000000000;
    #10 assign a = 64'h0007FFFFFFFFFFFF; assign b = 64'h400FFFFFFFFFFFFF;

    #10 $display("\n2**-1023 * 2**0:");
    #10 assign a = 64'h0008000000000000; assign b = 64'h3FF0000000000000;
    #10 assign a = 64'h000FFFFFFFFFFFFF; assign b = 64'h3FFFFFFFFFFFFFFF;

    #10 $display("\n2**-1022 * 2**-1:");
    #10 assign a = 64'h0010000000000000; assign b = 64'h3FE0000000000000;
    #10 assign a = 64'h001FFFFFFFFFFFFF; assign b = 64'h3FEFFFFFFFFFFFFF;

    #10 $display("\n2**-1021 * 2**-2:");
    #10 assign a = 64'h0020000000000000; assign b = 64'h3FD0000000000000;
    #10 assign a = 64'h002FFFFFFFFFFFFF; assign b = 64'h3FDFFFFFFFFFFFFF;

    #10 $display("\n2**-1020 * 2**-3:");
    #10 assign a = 64'h0030000000000000; assign b = 64'h3FC0000000000000;
    #10 assign a = 64'h003FFFFFFFFFFFFF; assign b = 64'h3FCFFFFFFFFFFFFF;

    #10 $display("\n2**-1019 * 2**-4:");
    #10 assign a = 64'h0040000000000000; assign b = 64'h3FB0000000000000;
    #10 assign a = 64'h004FFFFFFFFFFFFF; assign b = 64'h3FBFFFFFFFFFFFFF;

    #10 $display("\n2**-1018 * 2**-5:");
    #10 assign a = 64'h0050000000000000; assign b = 64'h3FA0000000000000;
    #10 assign a = 64'h005FFFFFFFFFFFFF; assign b = 64'h3FAFFFFFFFFFFFFF;

    #10 $display("\n2**-1017 * 2**-6:");
    #10 assign a = 64'h0060000000000000; assign b = 64'h3F90000000000000;
    #10 assign a = 64'h006FFFFFFFFFFFFF; assign b = 64'h3F9FFFFFFFFFFFFF;

    #10 $display("\n2**-1016 * 2**-7:");
    #10 assign a = 64'h0070000000000000; assign b = 64'h3F80000000000000;
    #10 assign a = 64'h007FFFFFFFFFFFFF; assign b = 64'h3F8FFFFFFFFFFFFF;

    #10 $display("\n2**-1015 * 2**-8:");
    #10 assign a = 64'h0080000000000000; assign b = 64'h3F70000000000000;
    #10 assign a = 64'h008FFFFFFFFFFFFF; assign b = 64'h3F7FFFFFFFFFFFFF;

    #10 $display("\n2**-1014 * 2**-9:");
    #10 assign a = 64'h0090000000000000; assign b = 64'h3F60000000000000;
    #10 assign a = 64'h009FFFFFFFFFFFFF; assign b = 64'h3F6FFFFFFFFFFFFF;

    #10 $display("\n2**-1013 * 2**-10:");
    #10 assign a = 64'h00A0000000000000; assign b = 64'h3F50000000000000;
    #10 assign a = 64'h00AFFFFFFFFFFFFF; assign b = 64'h3F5FFFFFFFFFFFFF;

    #10 $display("\n2**-1012 * 2**-11:");
    #10 assign a = 64'h00B0000000000000; assign b = 64'h3F40000000000000;
    #10 assign a = 64'h00BFFFFFFFFFFFFF; assign b = 64'h3F4FFFFFFFFFFFFF;

    #10 $display("\n2**-1011 * 2**-12:");
    #10 assign a = 64'h00C0000000000000; assign b = 64'h3F30000000000000;
    #10 assign a = 64'h00CFFFFFFFFFFFFF; assign b = 64'h3F3FFFFFFFFFFFFF;

    #10 $display("\n2**-1010 * 2**-13:");
    #10 assign a = 64'h00D0000000000000; assign b = 64'h3F20000000000000;
    #10 assign a = 64'h00DFFFFFFFFFFFFF; assign b = 64'h3F2FFFFFFFFFFFFF;

    #10 $display("\n2**-1009 * 2**-14:");
    #10 assign a = 64'h00E0000000000000; assign b = 64'h3F10000000000000;
    #10 assign a = 64'h00EFFFFFFFFFFFFF; assign b = 64'h3F1FFFFFFFFFFFFF;

    #10 $display("\n2**-1008 * 2**-15:");
    #10 assign a = 64'h00F0000000000000; assign b = 64'h3F00000000000000;
    #10 assign a = 64'h00FFFFFFFFFFFFFF; assign b = 64'h3F0FFFFFFFFFFFFF;

    #10 $display("\n2**-1007 * 2**-16:");
    #10 assign a = 64'h0100000000000000; assign b = 64'h3EF0000000000000;
    #10 assign a = 64'h010FFFFFFFFFFFFF; assign b = 64'h3EFFFFFFFFFFFFFF;

    #10 $display("\n2**-1006 * 2**-17:");
    #10 assign a = 64'h0110000000000000; assign b = 64'h3EE0000000000000;
    #10 assign a = 64'h011FFFFFFFFFFFFF; assign b = 64'h3EEFFFFFFFFFFFFF;

    #10 $display("\n2**-1005 * 2**-18:");
    #10 assign a = 64'h0120000000000000; assign b = 64'h3ED0000000000000;
    #10 assign a = 64'h012FFFFFFFFFFFFF; assign b = 64'h3EDFFFFFFFFFFFFF;

    #10 $display("\n2**-1004 * 2**-19:");
    #10 assign a = 64'h0130000000000000; assign b = 64'h3EC0000000000000;
    #10 assign a = 64'h013FFFFFFFFFFFFF; assign b = 64'h3ECFFFFFFFFFFFFF;

    #10 $display("\n2**-1003 * 2**-20:");
    #10 assign a = 64'h0140000000000000; assign b = 64'h3EB0000000000000;
    #10 assign a = 64'h014FFFFFFFFFFFFF; assign b = 64'h3EBFFFFFFFFFFFFF;

    #10 $display("\n2**-1002 * 2**-21:");
    #10 assign a = 64'h0150000000000000; assign b = 64'h3EA0000000000000;
    #10 assign a = 64'h015FFFFFFFFFFFFF; assign b = 64'h3EAFFFFFFFFFFFFF;

    #10 $display("\n2**-1001 * 2**-22:");
    #10 assign a = 64'h0160000000000000; assign b = 64'h3E90000000000000;
    #10 assign a = 64'h016FFFFFFFFFFFFF; assign b = 64'h3E9FFFFFFFFFFFFF;

    #10 $display("\n2**-1000 * 2**-23:");
    #10 assign a = 64'h0170000000000000; assign b = 64'h3E80000000000000;
    #10 assign a = 64'h017FFFFFFFFFFFFF; assign b = 64'h3E8FFFFFFFFFFFFF;

    #10 $display("\n2**-999 * 2**-24:");
    #10 assign a = 64'h0180000000000000; assign b = 64'h3E70000000000000;
    #10 assign a = 64'h018FFFFFFFFFFFFF; assign b = 64'h3E7FFFFFFFFFFFFF;

    #10 $display("\n2**-998 * 2**-25:");
    #10 assign a = 64'h0190000000000000; assign b = 64'h3E60000000000000;
    #10 assign a = 64'h019FFFFFFFFFFFFF; assign b = 64'h3E6FFFFFFFFFFFFF;

    #10 $display("\n2**-997 * 2**-26:");
    #10 assign a = 64'h01A0000000000000; assign b = 64'h3E50000000000000;
    #10 assign a = 64'h01AFFFFFFFFFFFFF; assign b = 64'h3E5FFFFFFFFFFFFF;

    #10 $display("\n2**-996 * 2**-27:");
    #10 assign a = 64'h01B0000000000000; assign b = 64'h3E40000000000000;
    #10 assign a = 64'h01BFFFFFFFFFFFFF; assign b = 64'h3E4FFFFFFFFFFFFF;

    #10 $display("\n2**-995 * 2**-28:");
    #10 assign a = 64'h01C0000000000000; assign b = 64'h3E30000000000000;
    #10 assign a = 64'h01CFFFFFFFFFFFFF; assign b = 64'h3E3FFFFFFFFFFFFF;

    #10 $display("\n2**-994 * 2**-29:");
    #10 assign a = 64'h01D0000000000000; assign b = 64'h3E20000000000000;
    #10 assign a = 64'h01DFFFFFFFFFFFFF; assign b = 64'h3E2FFFFFFFFFFFFF;

    #10 $display("\n2**-993 * 2**-30:");
    #10 assign a = 64'h01E0000000000000; assign b = 64'h3E10000000000000;
    #10 assign a = 64'h01EFFFFFFFFFFFFF; assign b = 64'h3E1FFFFFFFFFFFFF;

    #10 $display("\n2**-992 * 2**-31:");
    #10 assign a = 64'h01F0000000000000; assign b = 64'h3E00000000000000;
    #10 assign a = 64'h01FFFFFFFFFFFFFF; assign b = 64'h3E0FFFFFFFFFFFFF;

    #10 $display("\n2**-991 * 2**-32:");
    #10 assign a = 64'h0200000000000000; assign b = 64'h3DF0000000000000;
    #10 assign a = 64'h020FFFFFFFFFFFFF; assign b = 64'h3DFFFFFFFFFFFFFF;

    #10 $display("\n2**-990 * 2**-33:");
    #10 assign a = 64'h0210000000000000; assign b = 64'h3DE0000000000000;
    #10 assign a = 64'h021FFFFFFFFFFFFF; assign b = 64'h3DEFFFFFFFFFFFFF;

    #10 $display("\n2**-989 * 2**-34:");
    #10 assign a = 64'h0220000000000000; assign b = 64'h3DD0000000000000;
    #10 assign a = 64'h022FFFFFFFFFFFFF; assign b = 64'h3DDFFFFFFFFFFFFF;

    #10 $display("\n2**-988 * 2**-35:");
    #10 assign a = 64'h0230000000000000; assign b = 64'h3DC0000000000000;
    #10 assign a = 64'h023FFFFFFFFFFFFF; assign b = 64'h3DCFFFFFFFFFFFFF;

    #10 $display("\n2**-987 * 2**-36:");
    #10 assign a = 64'h0240000000000000; assign b = 64'h3DB0000000000000;
    #10 assign a = 64'h024FFFFFFFFFFFFF; assign b = 64'h3DBFFFFFFFFFFFFF;

    #10 $display("\n2**-986 * 2**-37:");
    #10 assign a = 64'h0250000000000000; assign b = 64'h3DA0000000000000;
    #10 assign a = 64'h025FFFFFFFFFFFFF; assign b = 64'h3DAFFFFFFFFFFFFF;

    #10 $display("\n2**-985 * 2**-38:");
    #10 assign a = 64'h0260000000000000; assign b = 64'h3D90000000000000;
    #10 assign a = 64'h026FFFFFFFFFFFFF; assign b = 64'h3D9FFFFFFFFFFFFF;

    #10 $display("\n2**-984 * 2**-39:");
    #10 assign a = 64'h0270000000000000; assign b = 64'h3D80000000000000;
    #10 assign a = 64'h027FFFFFFFFFFFFF; assign b = 64'h3D8FFFFFFFFFFFFF;

    #10 $display("\n2**-983 * 2**-40:");
    #10 assign a = 64'h0280000000000000; assign b = 64'h3D70000000000000;
    #10 assign a = 64'h028FFFFFFFFFFFFF; assign b = 64'h3D7FFFFFFFFFFFFF;

    #10 $display("\n2**-982 * 2**-41:");
    #10 assign a = 64'h0290000000000000; assign b = 64'h3D60000000000000;
    #10 assign a = 64'h029FFFFFFFFFFFFF; assign b = 64'h3D6FFFFFFFFFFFFF;

    #10 $display("\n2**-981 * 2**-42:");
    #10 assign a = 64'h02A0000000000000; assign b = 64'h3D50000000000000;
    #10 assign a = 64'h02AFFFFFFFFFFFFF; assign b = 64'h3D5FFFFFFFFFFFFF;

    #10 $display("\n2**-980 * 2**-43:");
    #10 assign a = 64'h02B0000000000000; assign b = 64'h3D40000000000000;
    #10 assign a = 64'h02BFFFFFFFFFFFFF; assign b = 64'h3D4FFFFFFFFFFFFF;

    #10 $display("\n2**-979 * 2**-44:");
    #10 assign a = 64'h02C0000000000000; assign b = 64'h3D30000000000000;
    #10 assign a = 64'h02CFFFFFFFFFFFFF; assign b = 64'h3D3FFFFFFFFFFFFF;

    #10 $display("\n2**-978 * 2**-45:");
    #10 assign a = 64'h02D0000000000000; assign b = 64'h3D20000000000000;
    #10 assign a = 64'h02DFFFFFFFFFFFFF; assign b = 64'h3D2FFFFFFFFFFFFF;

    #10 $display("\n2**-977 * 2**-46:");
    #10 assign a = 64'h02E0000000000000; assign b = 64'h3D10000000000000;
    #10 assign a = 64'h02EFFFFFFFFFFFFF; assign b = 64'h3D1FFFFFFFFFFFFF;

    #10 $display("\n2**-976 * 2**-47:");
    #10 assign a = 64'h02F0000000000000; assign b = 64'h3D00000000000000;
    #10 assign a = 64'h02FFFFFFFFFFFFFF; assign b = 64'h3D0FFFFFFFFFFFFF;

    #10 $display("\n2**-975 * 2**-48:");
    #10 assign a = 64'h0300000000000000; assign b = 64'h3CF0000000000000;
    #10 assign a = 64'h030FFFFFFFFFFFFF; assign b = 64'h3CFFFFFFFFFFFFFF;

    #10 $display("\n2**-974 * 2**-49:");
    #10 assign a = 64'h0310000000000000; assign b = 64'h3CE0000000000000;
    #10 assign a = 64'h031FFFFFFFFFFFFF; assign b = 64'h3CEFFFFFFFFFFFFF;

    #10 $display("\n2**-973 * 2**-50:");
    #10 assign a = 64'h0320000000000000; assign b = 64'h3CD0000000000000;
    #10 assign a = 64'h032FFFFFFFFFFFFF; assign b = 64'h3CDFFFFFFFFFFFFF;

    #10 $display("\n2**-972 * 2**-51:");
    #10 assign a = 64'h0330000000000000; assign b = 64'h3CC0000000000000;
    #10 assign a = 64'h033FFFFFFFFFFFFF; assign b = 64'h3CCFFFFFFFFFFFFF;

    #10 $display("\n2**-971 * 2**-52:");
    #10 assign a = 64'h0340000000000000; assign b = 64'h3CB0000000000000;
    #10 assign a = 64'h034FFFFFFFFFFFFF; assign b = 64'h3CBFFFFFFFFFFFFF;

    #10 $display("\n2**-970 * 2**-53:");
    #10 assign a = 64'h0350000000000000; assign b = 64'h3CA0000000000000;
    #10 assign a = 64'h035FFFFFFFFFFFFF; assign b = 64'h3CAFFFFFFFFFFFFF;

    #10 $display("\n2**-969 * 2**-54:");
    #10 assign a = 64'h0360000000000000; assign b = 64'h3C90000000000000;
    #10 assign a = 64'h036FFFFFFFFFFFFF; assign b = 64'h3C9FFFFFFFFFFFFF;

    #10 $display("\n2**-968 * 2**-55:");
    #10 assign a = 64'h0370000000000000; assign b = 64'h3C80000000000000;
    #10 assign a = 64'h037FFFFFFFFFFFFF; assign b = 64'h3C8FFFFFFFFFFFFF;

    #10 $display("\n2**-967 * 2**-56:");
    #10 assign a = 64'h0380000000000000; assign b = 64'h3C70000000000000;
    #10 assign a = 64'h038FFFFFFFFFFFFF; assign b = 64'h3C7FFFFFFFFFFFFF;

    #10 $display("\n2**-966 * 2**-57:");
    #10 assign a = 64'h0390000000000000; assign b = 64'h3C60000000000000;
    #10 assign a = 64'h039FFFFFFFFFFFFF; assign b = 64'h3C6FFFFFFFFFFFFF;

    #10 $display("\n2**-965 * 2**-58:");
    #10 assign a = 64'h03A0000000000000; assign b = 64'h3C50000000000000;
    #10 assign a = 64'h03AFFFFFFFFFFFFF; assign b = 64'h3C5FFFFFFFFFFFFF;

    #10 $display("\n2**-964 * 2**-59:");
    #10 assign a = 64'h03B0000000000000; assign b = 64'h3C40000000000000;
    #10 assign a = 64'h03BFFFFFFFFFFFFF; assign b = 64'h3C4FFFFFFFFFFFFF;

    #10 $display("\n2**-963 * 2**-60:");
    #10 assign a = 64'h03C0000000000000; assign b = 64'h3C30000000000000;
    #10 assign a = 64'h03CFFFFFFFFFFFFF; assign b = 64'h3C3FFFFFFFFFFFFF;

    #10 $display("\n2**-962 * 2**-61:");
    #10 assign a = 64'h03D0000000000000; assign b = 64'h3C20000000000000;
    #10 assign a = 64'h03DFFFFFFFFFFFFF; assign b = 64'h3C2FFFFFFFFFFFFF;

    #10 $display("\n2**-961 * 2**-62:");
    #10 assign a = 64'h03E0000000000000; assign b = 64'h3C10000000000000;
    #10 assign a = 64'h03EFFFFFFFFFFFFF; assign b = 64'h3C1FFFFFFFFFFFFF;

    #10 $display("\n2**-960 * 2**-63:");
    #10 assign a = 64'h03F0000000000000; assign b = 64'h3C00000000000000;
    #10 assign a = 64'h03FFFFFFFFFFFFFF; assign b = 64'h3C0FFFFFFFFFFFFF;

    #10 $display("\n2**-959 * 2**-64:");
    #10 assign a = 64'h0400000000000000; assign b = 64'h3BF0000000000000;
    #10 assign a = 64'h040FFFFFFFFFFFFF; assign b = 64'h3BFFFFFFFFFFFFFF;

    #10 $display("\n2**-958 * 2**-65:");
    #10 assign a = 64'h0410000000000000; assign b = 64'h3BE0000000000000;
    #10 assign a = 64'h041FFFFFFFFFFFFF; assign b = 64'h3BEFFFFFFFFFFFFF;

    #10 $display("\n2**-957 * 2**-66:");
    #10 assign a = 64'h0420000000000000; assign b = 64'h3BD0000000000000;
    #10 assign a = 64'h042FFFFFFFFFFFFF; assign b = 64'h3BDFFFFFFFFFFFFF;

    #10 $display("\n2**-956 * 2**-67:");
    #10 assign a = 64'h0430000000000000; assign b = 64'h3BC0000000000000;
    #10 assign a = 64'h043FFFFFFFFFFFFF; assign b = 64'h3BCFFFFFFFFFFFFF;

    #10 $display("\n2**-955 * 2**-68:");
    #10 assign a = 64'h0440000000000000; assign b = 64'h3BB0000000000000;
    #10 assign a = 64'h044FFFFFFFFFFFFF; assign b = 64'h3BBFFFFFFFFFFFFF;

    #10 $display("\n2**-954 * 2**-69:");
    #10 assign a = 64'h0450000000000000; assign b = 64'h3BA0000000000000;
    #10 assign a = 64'h045FFFFFFFFFFFFF; assign b = 64'h3BAFFFFFFFFFFFFF;

    #10 $display("\n2**-953 * 2**-70:");
    #10 assign a = 64'h0460000000000000; assign b = 64'h3B90000000000000;
    #10 assign a = 64'h046FFFFFFFFFFFFF; assign b = 64'h3B9FFFFFFFFFFFFF;

    #10 $display("\n2**-952 * 2**-71:");
    #10 assign a = 64'h0470000000000000; assign b = 64'h3B80000000000000;
    #10 assign a = 64'h047FFFFFFFFFFFFF; assign b = 64'h3B8FFFFFFFFFFFFF;

    #10 $display("\n2**-951 * 2**-72:");
    #10 assign a = 64'h0480000000000000; assign b = 64'h3B70000000000000;
    #10 assign a = 64'h048FFFFFFFFFFFFF; assign b = 64'h3B7FFFFFFFFFFFFF;

    #10 $display("\n2**-950 * 2**-73:");
    #10 assign a = 64'h0490000000000000; assign b = 64'h3B60000000000000;
    #10 assign a = 64'h049FFFFFFFFFFFFF; assign b = 64'h3B6FFFFFFFFFFFFF;

    #10 $display("\n2**-949 * 2**-74:");
    #10 assign a = 64'h04A0000000000000; assign b = 64'h3B50000000000000;
    #10 assign a = 64'h04AFFFFFFFFFFFFF; assign b = 64'h3B5FFFFFFFFFFFFF;

    #10 $display("\n2**-948 * 2**-75:");
    #10 assign a = 64'h04B0000000000000; assign b = 64'h3B40000000000000;
    #10 assign a = 64'h04BFFFFFFFFFFFFF; assign b = 64'h3B4FFFFFFFFFFFFF;

    #10 $display("\n2**-947 * 2**-76:");
    #10 assign a = 64'h04C0000000000000; assign b = 64'h3B30000000000000;
    #10 assign a = 64'h04CFFFFFFFFFFFFF; assign b = 64'h3B3FFFFFFFFFFFFF;

    #10 $display("\n2**-946 * 2**-77:");
    #10 assign a = 64'h04D0000000000000; assign b = 64'h3B20000000000000;
    #10 assign a = 64'h04DFFFFFFFFFFFFF; assign b = 64'h3B2FFFFFFFFFFFFF;

    #10 $display("\n2**-945 * 2**-78:");
    #10 assign a = 64'h04E0000000000000; assign b = 64'h3B10000000000000;
    #10 assign a = 64'h04EFFFFFFFFFFFFF; assign b = 64'h3B1FFFFFFFFFFFFF;

    #10 $display("\n2**-944 * 2**-79:");
    #10 assign a = 64'h04F0000000000000; assign b = 64'h3B00000000000000;
    #10 assign a = 64'h04FFFFFFFFFFFFFF; assign b = 64'h3B0FFFFFFFFFFFFF;

    #10 $display("\n2**-943 * 2**-80:");
    #10 assign a = 64'h0500000000000000; assign b = 64'h3AF0000000000000;
    #10 assign a = 64'h050FFFFFFFFFFFFF; assign b = 64'h3AFFFFFFFFFFFFFF;

    #10 $display("\n2**-942 * 2**-81:");
    #10 assign a = 64'h0510000000000000; assign b = 64'h3AE0000000000000;
    #10 assign a = 64'h051FFFFFFFFFFFFF; assign b = 64'h3AEFFFFFFFFFFFFF;

    #10 $display("\n2**-941 * 2**-82:");
    #10 assign a = 64'h0520000000000000; assign b = 64'h3AD0000000000000;
    #10 assign a = 64'h052FFFFFFFFFFFFF; assign b = 64'h3ADFFFFFFFFFFFFF;

    #10 $display("\n2**-940 * 2**-83:");
    #10 assign a = 64'h0530000000000000; assign b = 64'h3AC0000000000000;
    #10 assign a = 64'h053FFFFFFFFFFFFF; assign b = 64'h3ACFFFFFFFFFFFFF;

    #10 $display("\n2**-939 * 2**-84:");
    #10 assign a = 64'h0540000000000000; assign b = 64'h3AB0000000000000;
    #10 assign a = 64'h054FFFFFFFFFFFFF; assign b = 64'h3ABFFFFFFFFFFFFF;

    #10 $display("\n2**-938 * 2**-85:");
    #10 assign a = 64'h0550000000000000; assign b = 64'h3AA0000000000000;
    #10 assign a = 64'h055FFFFFFFFFFFFF; assign b = 64'h3AAFFFFFFFFFFFFF;

    #10 $display("\n2**-937 * 2**-86:");
    #10 assign a = 64'h0560000000000000; assign b = 64'h3A90000000000000;
    #10 assign a = 64'h056FFFFFFFFFFFFF; assign b = 64'h3A9FFFFFFFFFFFFF;

    #10 $display("\n2**-936 * 2**-87:");
    #10 assign a = 64'h0570000000000000; assign b = 64'h3A80000000000000;
    #10 assign a = 64'h057FFFFFFFFFFFFF; assign b = 64'h3A8FFFFFFFFFFFFF;

    #10 $display("\n2**-935 * 2**-88:");
    #10 assign a = 64'h0580000000000000; assign b = 64'h3A70000000000000;
    #10 assign a = 64'h058FFFFFFFFFFFFF; assign b = 64'h3A7FFFFFFFFFFFFF;

    #10 $display("\n2**-934 * 2**-89:");
    #10 assign a = 64'h0590000000000000; assign b = 64'h3A60000000000000;
    #10 assign a = 64'h059FFFFFFFFFFFFF; assign b = 64'h3A6FFFFFFFFFFFFF;

    #10 $display("\n2**-933 * 2**-90:");
    #10 assign a = 64'h05A0000000000000; assign b = 64'h3A50000000000000;
    #10 assign a = 64'h05AFFFFFFFFFFFFF; assign b = 64'h3A5FFFFFFFFFFFFF;

    #10 $display("\n2**-932 * 2**-91:");
    #10 assign a = 64'h05B0000000000000; assign b = 64'h3A40000000000000;
    #10 assign a = 64'h05BFFFFFFFFFFFFF; assign b = 64'h3A4FFFFFFFFFFFFF;

    #10 $display("\n2**-931 * 2**-92:");
    #10 assign a = 64'h05C0000000000000; assign b = 64'h3A30000000000000;
    #10 assign a = 64'h05CFFFFFFFFFFFFF; assign b = 64'h3A3FFFFFFFFFFFFF;

    #10 $display("\n2**-930 * 2**-93:");
    #10 assign a = 64'h05D0000000000000; assign b = 64'h3A20000000000000;
    #10 assign a = 64'h05DFFFFFFFFFFFFF; assign b = 64'h3A2FFFFFFFFFFFFF;

    #10 $display("\n2**-929 * 2**-94:");
    #10 assign a = 64'h05E0000000000000; assign b = 64'h3A10000000000000;
    #10 assign a = 64'h05EFFFFFFFFFFFFF; assign b = 64'h3A1FFFFFFFFFFFFF;

    #10 $display("\n2**-928 * 2**-95:");
    #10 assign a = 64'h05F0000000000000; assign b = 64'h3A00000000000000;
    #10 assign a = 64'h05FFFFFFFFFFFFFF; assign b = 64'h3A0FFFFFFFFFFFFF;

    #10 $display("\n2**-927 * 2**-96:");
    #10 assign a = 64'h0600000000000000; assign b = 64'h39F0000000000000;
    #10 assign a = 64'h060FFFFFFFFFFFFF; assign b = 64'h39FFFFFFFFFFFFFF;

    #10 $display("\n2**-926 * 2**-97:");
    #10 assign a = 64'h0610000000000000; assign b = 64'h39E0000000000000;
    #10 assign a = 64'h061FFFFFFFFFFFFF; assign b = 64'h39EFFFFFFFFFFFFF;

    #10 $display("\n2**-925 * 2**-98:");
    #10 assign a = 64'h0620000000000000; assign b = 64'h39D0000000000000;
    #10 assign a = 64'h062FFFFFFFFFFFFF; assign b = 64'h39DFFFFFFFFFFFFF;

    #10 $display("\n2**-924 * 2**-99:");
    #10 assign a = 64'h0630000000000000; assign b = 64'h39C0000000000000;
    #10 assign a = 64'h063FFFFFFFFFFFFF; assign b = 64'h39CFFFFFFFFFFFFF;

    #10 $display("\n2**-923 * 2**-100:");
    #10 assign a = 64'h0640000000000000; assign b = 64'h39B0000000000000;
    #10 assign a = 64'h064FFFFFFFFFFFFF; assign b = 64'h39BFFFFFFFFFFFFF;

    #10 $display("\n2**-922 * 2**-101:");
    #10 assign a = 64'h0650000000000000; assign b = 64'h39A0000000000000;
    #10 assign a = 64'h065FFFFFFFFFFFFF; assign b = 64'h39AFFFFFFFFFFFFF;

    #10 $display("\n2**-921 * 2**-102:");
    #10 assign a = 64'h0660000000000000; assign b = 64'h3990000000000000;
    #10 assign a = 64'h066FFFFFFFFFFFFF; assign b = 64'h399FFFFFFFFFFFFF;

    #10 $display("\n2**-920 * 2**-103:");
    #10 assign a = 64'h0670000000000000; assign b = 64'h3980000000000000;
    #10 assign a = 64'h067FFFFFFFFFFFFF; assign b = 64'h398FFFFFFFFFFFFF;

    #10 $display("\n2**-919 * 2**-104:");
    #10 assign a = 64'h0680000000000000; assign b = 64'h3970000000000000;
    #10 assign a = 64'h068FFFFFFFFFFFFF; assign b = 64'h397FFFFFFFFFFFFF;

    #10 $display("\n2**-918 * 2**-105:");
    #10 assign a = 64'h0690000000000000; assign b = 64'h3960000000000000;
    #10 assign a = 64'h069FFFFFFFFFFFFF; assign b = 64'h396FFFFFFFFFFFFF;

    #10 $display("\n2**-917 * 2**-106:");
    #10 assign a = 64'h06A0000000000000; assign b = 64'h3950000000000000;
    #10 assign a = 64'h06AFFFFFFFFFFFFF; assign b = 64'h395FFFFFFFFFFFFF;

    #10 $display("\n2**-916 * 2**-107:");
    #10 assign a = 64'h06B0000000000000; assign b = 64'h3940000000000000;
    #10 assign a = 64'h06BFFFFFFFFFFFFF; assign b = 64'h394FFFFFFFFFFFFF;

    #10 $display("\n2**-915 * 2**-108:");
    #10 assign a = 64'h06C0000000000000; assign b = 64'h3930000000000000;
    #10 assign a = 64'h06CFFFFFFFFFFFFF; assign b = 64'h393FFFFFFFFFFFFF;

    #10 $display("\n2**-914 * 2**-109:");
    #10 assign a = 64'h06D0000000000000; assign b = 64'h3920000000000000;
    #10 assign a = 64'h06DFFFFFFFFFFFFF; assign b = 64'h392FFFFFFFFFFFFF;

    #10 $display("\n2**-913 * 2**-110:");
    #10 assign a = 64'h06E0000000000000; assign b = 64'h3910000000000000;
    #10 assign a = 64'h06EFFFFFFFFFFFFF; assign b = 64'h391FFFFFFFFFFFFF;

    #10 $display("\n2**-912 * 2**-111:");
    #10 assign a = 64'h06F0000000000000; assign b = 64'h3900000000000000;
    #10 assign a = 64'h06FFFFFFFFFFFFFF; assign b = 64'h390FFFFFFFFFFFFF;

    #10 $display("\n2**-911 * 2**-112:");
    #10 assign a = 64'h0700000000000000; assign b = 64'h38F0000000000000;
    #10 assign a = 64'h070FFFFFFFFFFFFF; assign b = 64'h38FFFFFFFFFFFFFF;

    #10 $display("\n2**-910 * 2**-113:");
    #10 assign a = 64'h0710000000000000; assign b = 64'h38E0000000000000;
    #10 assign a = 64'h071FFFFFFFFFFFFF; assign b = 64'h38EFFFFFFFFFFFFF;

    #10 $display("\n2**-909 * 2**-114:");
    #10 assign a = 64'h0720000000000000; assign b = 64'h38D0000000000000;
    #10 assign a = 64'h072FFFFFFFFFFFFF; assign b = 64'h38DFFFFFFFFFFFFF;

    #10 $display("\n2**-908 * 2**-115:");
    #10 assign a = 64'h0730000000000000; assign b = 64'h38C0000000000000;
    #10 assign a = 64'h073FFFFFFFFFFFFF; assign b = 64'h38CFFFFFFFFFFFFF;

    #10 $display("\n2**-907 * 2**-116:");
    #10 assign a = 64'h0740000000000000; assign b = 64'h38B0000000000000;
    #10 assign a = 64'h074FFFFFFFFFFFFF; assign b = 64'h38BFFFFFFFFFFFFF;

    #10 $display("\n2**-906 * 2**-117:");
    #10 assign a = 64'h0750000000000000; assign b = 64'h38A0000000000000;
    #10 assign a = 64'h075FFFFFFFFFFFFF; assign b = 64'h38AFFFFFFFFFFFFF;

    #10 $display("\n2**-905 * 2**-118:");
    #10 assign a = 64'h0760000000000000; assign b = 64'h3890000000000000;
    #10 assign a = 64'h076FFFFFFFFFFFFF; assign b = 64'h389FFFFFFFFFFFFF;

    #10 $display("\n2**-904 * 2**-119:");
    #10 assign a = 64'h0770000000000000; assign b = 64'h3880000000000000;
    #10 assign a = 64'h077FFFFFFFFFFFFF; assign b = 64'h388FFFFFFFFFFFFF;

    #10 $display("\n2**-903 * 2**-120:");
    #10 assign a = 64'h0780000000000000; assign b = 64'h3870000000000000;
    #10 assign a = 64'h078FFFFFFFFFFFFF; assign b = 64'h387FFFFFFFFFFFFF;

    #10 $display("\n2**-902 * 2**-121:");
    #10 assign a = 64'h0790000000000000; assign b = 64'h3860000000000000;
    #10 assign a = 64'h079FFFFFFFFFFFFF; assign b = 64'h386FFFFFFFFFFFFF;

    #10 $display("\n2**-901 * 2**-122:");
    #10 assign a = 64'h07A0000000000000; assign b = 64'h3850000000000000;
    #10 assign a = 64'h07AFFFFFFFFFFFFF; assign b = 64'h385FFFFFFFFFFFFF;

    #10 $display("\n2**-900 * 2**-123:");
    #10 assign a = 64'h07B0000000000000; assign b = 64'h3840000000000000;
    #10 assign a = 64'h07BFFFFFFFFFFFFF; assign b = 64'h384FFFFFFFFFFFFF;

    #10 $display("\n2**-899 * 2**-124:");
    #10 assign a = 64'h07C0000000000000; assign b = 64'h3830000000000000;
    #10 assign a = 64'h07CFFFFFFFFFFFFF; assign b = 64'h383FFFFFFFFFFFFF;

    #10 $display("\n2**-898 * 2**-125:");
    #10 assign a = 64'h07D0000000000000; assign b = 64'h3820000000000000;
    #10 assign a = 64'h07DFFFFFFFFFFFFF; assign b = 64'h382FFFFFFFFFFFFF;

    #10 $display("\n2**-897 * 2**-126:");
    #10 assign a = 64'h07E0000000000000; assign b = 64'h3810000000000000;
    #10 assign a = 64'h07EFFFFFFFFFFFFF; assign b = 64'h381FFFFFFFFFFFFF;

    #10 $display("\n2**-896 * 2**-127:");
    #10 assign a = 64'h07F0000000000000; assign b = 64'h3800000000000000;
    #10 assign a = 64'h07FFFFFFFFFFFFFF; assign b = 64'h380FFFFFFFFFFFFF;

    #10 $display("\n2**-895 * 2**-128:");
    #10 assign a = 64'h0800000000000000; assign b = 64'h37F0000000000000;
    #10 assign a = 64'h080FFFFFFFFFFFFF; assign b = 64'h37FFFFFFFFFFFFFF;

    #10 $display("\n2**-894 * 2**-129:");
    #10 assign a = 64'h0810000000000000; assign b = 64'h37E0000000000000;
    #10 assign a = 64'h081FFFFFFFFFFFFF; assign b = 64'h37EFFFFFFFFFFFFF;

    #10 $display("\n2**-893 * 2**-130:");
    #10 assign a = 64'h0820000000000000; assign b = 64'h37D0000000000000;
    #10 assign a = 64'h082FFFFFFFFFFFFF; assign b = 64'h37DFFFFFFFFFFFFF;

    #10 $display("\n2**-892 * 2**-131:");
    #10 assign a = 64'h0830000000000000; assign b = 64'h37C0000000000000;
    #10 assign a = 64'h083FFFFFFFFFFFFF; assign b = 64'h37CFFFFFFFFFFFFF;

    #10 $display("\n2**-891 * 2**-132:");
    #10 assign a = 64'h0840000000000000; assign b = 64'h37B0000000000000;
    #10 assign a = 64'h084FFFFFFFFFFFFF; assign b = 64'h37BFFFFFFFFFFFFF;

    #10 $display("\n2**-890 * 2**-133:");
    #10 assign a = 64'h0850000000000000; assign b = 64'h37A0000000000000;
    #10 assign a = 64'h085FFFFFFFFFFFFF; assign b = 64'h37AFFFFFFFFFFFFF;

    #10 $display("\n2**-889 * 2**-134:");
    #10 assign a = 64'h0860000000000000; assign b = 64'h3790000000000000;
    #10 assign a = 64'h086FFFFFFFFFFFFF; assign b = 64'h379FFFFFFFFFFFFF;

    #10 $display("\n2**-888 * 2**-135:");
    #10 assign a = 64'h0870000000000000; assign b = 64'h3780000000000000;
    #10 assign a = 64'h087FFFFFFFFFFFFF; assign b = 64'h378FFFFFFFFFFFFF;

    #10 $display("\n2**-887 * 2**-136:");
    #10 assign a = 64'h0880000000000000; assign b = 64'h3770000000000000;
    #10 assign a = 64'h088FFFFFFFFFFFFF; assign b = 64'h377FFFFFFFFFFFFF;

    #10 $display("\n2**-886 * 2**-137:");
    #10 assign a = 64'h0890000000000000; assign b = 64'h3760000000000000;
    #10 assign a = 64'h089FFFFFFFFFFFFF; assign b = 64'h376FFFFFFFFFFFFF;

    #10 $display("\n2**-885 * 2**-138:");
    #10 assign a = 64'h08A0000000000000; assign b = 64'h3750000000000000;
    #10 assign a = 64'h08AFFFFFFFFFFFFF; assign b = 64'h375FFFFFFFFFFFFF;

    #10 $display("\n2**-884 * 2**-139:");
    #10 assign a = 64'h08B0000000000000; assign b = 64'h3740000000000000;
    #10 assign a = 64'h08BFFFFFFFFFFFFF; assign b = 64'h374FFFFFFFFFFFFF;

    #10 $display("\n2**-883 * 2**-140:");
    #10 assign a = 64'h08C0000000000000; assign b = 64'h3730000000000000;
    #10 assign a = 64'h08CFFFFFFFFFFFFF; assign b = 64'h373FFFFFFFFFFFFF;

    #10 $display("\n2**-882 * 2**-141:");
    #10 assign a = 64'h08D0000000000000; assign b = 64'h3720000000000000;
    #10 assign a = 64'h08DFFFFFFFFFFFFF; assign b = 64'h372FFFFFFFFFFFFF;

    #10 $display("\n2**-881 * 2**-142:");
    #10 assign a = 64'h08E0000000000000; assign b = 64'h3710000000000000;
    #10 assign a = 64'h08EFFFFFFFFFFFFF; assign b = 64'h371FFFFFFFFFFFFF;

    #10 $display("\n2**-880 * 2**-143:");
    #10 assign a = 64'h08F0000000000000; assign b = 64'h3700000000000000;
    #10 assign a = 64'h08FFFFFFFFFFFFFF; assign b = 64'h370FFFFFFFFFFFFF;

    #10 $display("\n2**-879 * 2**-144:");
    #10 assign a = 64'h0900000000000000; assign b = 64'h36F0000000000000;
    #10 assign a = 64'h090FFFFFFFFFFFFF; assign b = 64'h36FFFFFFFFFFFFFF;

    #10 $display("\n2**-878 * 2**-145:");
    #10 assign a = 64'h0910000000000000; assign b = 64'h36E0000000000000;
    #10 assign a = 64'h091FFFFFFFFFFFFF; assign b = 64'h36EFFFFFFFFFFFFF;

    #10 $display("\n2**-877 * 2**-146:");
    #10 assign a = 64'h0920000000000000; assign b = 64'h36D0000000000000;
    #10 assign a = 64'h092FFFFFFFFFFFFF; assign b = 64'h36DFFFFFFFFFFFFF;

    #10 $display("\n2**-876 * 2**-147:");
    #10 assign a = 64'h0930000000000000; assign b = 64'h36C0000000000000;
    #10 assign a = 64'h093FFFFFFFFFFFFF; assign b = 64'h36CFFFFFFFFFFFFF;

    #10 $display("\n2**-875 * 2**-148:");
    #10 assign a = 64'h0940000000000000; assign b = 64'h36B0000000000000;
    #10 assign a = 64'h094FFFFFFFFFFFFF; assign b = 64'h36BFFFFFFFFFFFFF;

    #10 $display("\n2**-874 * 2**-149:");
    #10 assign a = 64'h0950000000000000; assign b = 64'h36A0000000000000;
    #10 assign a = 64'h095FFFFFFFFFFFFF; assign b = 64'h36AFFFFFFFFFFFFF;

    #10 $display("\n2**-873 * 2**-150:");
    #10 assign a = 64'h0960000000000000; assign b = 64'h3690000000000000;
    #10 assign a = 64'h096FFFFFFFFFFFFF; assign b = 64'h369FFFFFFFFFFFFF;

    #10 $display("\n2**-872 * 2**-151:");
    #10 assign a = 64'h0970000000000000; assign b = 64'h3680000000000000;
    #10 assign a = 64'h097FFFFFFFFFFFFF; assign b = 64'h368FFFFFFFFFFFFF;

    #10 $display("\n2**-871 * 2**-152:");
    #10 assign a = 64'h0980000000000000; assign b = 64'h3670000000000000;
    #10 assign a = 64'h098FFFFFFFFFFFFF; assign b = 64'h367FFFFFFFFFFFFF;

    #10 $display("\n2**-870 * 2**-153:");
    #10 assign a = 64'h0990000000000000; assign b = 64'h3660000000000000;
    #10 assign a = 64'h099FFFFFFFFFFFFF; assign b = 64'h366FFFFFFFFFFFFF;

    #10 $display("\n2**-869 * 2**-154:");
    #10 assign a = 64'h09A0000000000000; assign b = 64'h3650000000000000;
    #10 assign a = 64'h09AFFFFFFFFFFFFF; assign b = 64'h365FFFFFFFFFFFFF;

    #10 $display("\n2**-868 * 2**-155:");
    #10 assign a = 64'h09B0000000000000; assign b = 64'h3640000000000000;
    #10 assign a = 64'h09BFFFFFFFFFFFFF; assign b = 64'h364FFFFFFFFFFFFF;

    #10 $display("\n2**-867 * 2**-156:");
    #10 assign a = 64'h09C0000000000000; assign b = 64'h3630000000000000;
    #10 assign a = 64'h09CFFFFFFFFFFFFF; assign b = 64'h363FFFFFFFFFFFFF;

    #10 $display("\n2**-866 * 2**-157:");
    #10 assign a = 64'h09D0000000000000; assign b = 64'h3620000000000000;
    #10 assign a = 64'h09DFFFFFFFFFFFFF; assign b = 64'h362FFFFFFFFFFFFF;

    #10 $display("\n2**-865 * 2**-158:");
    #10 assign a = 64'h09E0000000000000; assign b = 64'h3610000000000000;
    #10 assign a = 64'h09EFFFFFFFFFFFFF; assign b = 64'h361FFFFFFFFFFFFF;

    #10 $display("\n2**-864 * 2**-159:");
    #10 assign a = 64'h09F0000000000000; assign b = 64'h3600000000000000;
    #10 assign a = 64'h09FFFFFFFFFFFFFF; assign b = 64'h360FFFFFFFFFFFFF;

    #10 $display("\n2**-863 * 2**-160:");
    #10 assign a = 64'h0A00000000000000; assign b = 64'h35F0000000000000;
    #10 assign a = 64'h0A0FFFFFFFFFFFFF; assign b = 64'h35FFFFFFFFFFFFFF;

    #10 $display("\n2**-862 * 2**-161:");
    #10 assign a = 64'h0A10000000000000; assign b = 64'h35E0000000000000;
    #10 assign a = 64'h0A1FFFFFFFFFFFFF; assign b = 64'h35EFFFFFFFFFFFFF;

    #10 $display("\n2**-861 * 2**-162:");
    #10 assign a = 64'h0A20000000000000; assign b = 64'h35D0000000000000;
    #10 assign a = 64'h0A2FFFFFFFFFFFFF; assign b = 64'h35DFFFFFFFFFFFFF;

    #10 $display("\n2**-860 * 2**-163:");
    #10 assign a = 64'h0A30000000000000; assign b = 64'h35C0000000000000;
    #10 assign a = 64'h0A3FFFFFFFFFFFFF; assign b = 64'h35CFFFFFFFFFFFFF;

    #10 $display("\n2**-859 * 2**-164:");
    #10 assign a = 64'h0A40000000000000; assign b = 64'h35B0000000000000;
    #10 assign a = 64'h0A4FFFFFFFFFFFFF; assign b = 64'h35BFFFFFFFFFFFFF;

    #10 $display("\n2**-858 * 2**-165:");
    #10 assign a = 64'h0A50000000000000; assign b = 64'h35A0000000000000;
    #10 assign a = 64'h0A5FFFFFFFFFFFFF; assign b = 64'h35AFFFFFFFFFFFFF;

    #10 $display("\n2**-857 * 2**-166:");
    #10 assign a = 64'h0A60000000000000; assign b = 64'h3590000000000000;
    #10 assign a = 64'h0A6FFFFFFFFFFFFF; assign b = 64'h359FFFFFFFFFFFFF;

    #10 $display("\n2**-856 * 2**-167:");
    #10 assign a = 64'h0A70000000000000; assign b = 64'h3580000000000000;
    #10 assign a = 64'h0A7FFFFFFFFFFFFF; assign b = 64'h358FFFFFFFFFFFFF;

    #10 $display("\n2**-855 * 2**-168:");
    #10 assign a = 64'h0A80000000000000; assign b = 64'h3570000000000000;
    #10 assign a = 64'h0A8FFFFFFFFFFFFF; assign b = 64'h357FFFFFFFFFFFFF;

    #10 $display("\n2**-854 * 2**-169:");
    #10 assign a = 64'h0A90000000000000; assign b = 64'h3560000000000000;
    #10 assign a = 64'h0A9FFFFFFFFFFFFF; assign b = 64'h356FFFFFFFFFFFFF;

    #10 $display("\n2**-853 * 2**-170:");
    #10 assign a = 64'h0AA0000000000000; assign b = 64'h3550000000000000;
    #10 assign a = 64'h0AAFFFFFFFFFFFFF; assign b = 64'h355FFFFFFFFFFFFF;

    #10 $display("\n2**-852 * 2**-171:");
    #10 assign a = 64'h0AB0000000000000; assign b = 64'h3540000000000000;
    #10 assign a = 64'h0ABFFFFFFFFFFFFF; assign b = 64'h354FFFFFFFFFFFFF;

    #10 $display("\n2**-851 * 2**-172:");
    #10 assign a = 64'h0AC0000000000000; assign b = 64'h3530000000000000;
    #10 assign a = 64'h0ACFFFFFFFFFFFFF; assign b = 64'h353FFFFFFFFFFFFF;

    #10 $display("\n2**-850 * 2**-173:");
    #10 assign a = 64'h0AD0000000000000; assign b = 64'h3520000000000000;
    #10 assign a = 64'h0ADFFFFFFFFFFFFF; assign b = 64'h352FFFFFFFFFFFFF;

    #10 $display("\n2**-849 * 2**-174:");
    #10 assign a = 64'h0AE0000000000000; assign b = 64'h3510000000000000;
    #10 assign a = 64'h0AEFFFFFFFFFFFFF; assign b = 64'h351FFFFFFFFFFFFF;

    #10 $display("\n2**-848 * 2**-175:");
    #10 assign a = 64'h0AF0000000000000; assign b = 64'h3500000000000000;
    #10 assign a = 64'h0AFFFFFFFFFFFFFF; assign b = 64'h350FFFFFFFFFFFFF;

    #10 $display("\n2**-847 * 2**-176:");
    #10 assign a = 64'h0B00000000000000; assign b = 64'h34F0000000000000;
    #10 assign a = 64'h0B0FFFFFFFFFFFFF; assign b = 64'h34FFFFFFFFFFFFFF;

    #10 $display("\n2**-846 * 2**-177:");
    #10 assign a = 64'h0B10000000000000; assign b = 64'h34E0000000000000;
    #10 assign a = 64'h0B1FFFFFFFFFFFFF; assign b = 64'h34EFFFFFFFFFFFFF;

    #10 $display("\n2**-845 * 2**-178:");
    #10 assign a = 64'h0B20000000000000; assign b = 64'h34D0000000000000;
    #10 assign a = 64'h0B2FFFFFFFFFFFFF; assign b = 64'h34DFFFFFFFFFFFFF;

    #10 $display("\n2**-844 * 2**-179:");
    #10 assign a = 64'h0B30000000000000; assign b = 64'h34C0000000000000;
    #10 assign a = 64'h0B3FFFFFFFFFFFFF; assign b = 64'h34CFFFFFFFFFFFFF;

    #10 $display("\n2**-843 * 2**-180:");
    #10 assign a = 64'h0B40000000000000; assign b = 64'h34B0000000000000;
    #10 assign a = 64'h0B4FFFFFFFFFFFFF; assign b = 64'h34BFFFFFFFFFFFFF;

    #10 $display("\n2**-842 * 2**-181:");
    #10 assign a = 64'h0B50000000000000; assign b = 64'h34A0000000000000;
    #10 assign a = 64'h0B5FFFFFFFFFFFFF; assign b = 64'h34AFFFFFFFFFFFFF;

    #10 $display("\n2**-841 * 2**-182:");
    #10 assign a = 64'h0B60000000000000; assign b = 64'h3490000000000000;
    #10 assign a = 64'h0B6FFFFFFFFFFFFF; assign b = 64'h349FFFFFFFFFFFFF;

    #10 $display("\n2**-840 * 2**-183:");
    #10 assign a = 64'h0B70000000000000; assign b = 64'h3480000000000000;
    #10 assign a = 64'h0B7FFFFFFFFFFFFF; assign b = 64'h348FFFFFFFFFFFFF;

    #10 $display("\n2**-839 * 2**-184:");
    #10 assign a = 64'h0B80000000000000; assign b = 64'h3470000000000000;
    #10 assign a = 64'h0B8FFFFFFFFFFFFF; assign b = 64'h347FFFFFFFFFFFFF;

    #10 $display("\n2**-838 * 2**-185:");
    #10 assign a = 64'h0B90000000000000; assign b = 64'h3460000000000000;
    #10 assign a = 64'h0B9FFFFFFFFFFFFF; assign b = 64'h346FFFFFFFFFFFFF;

    #10 $display("\n2**-837 * 2**-186:");
    #10 assign a = 64'h0BA0000000000000; assign b = 64'h3450000000000000;
    #10 assign a = 64'h0BAFFFFFFFFFFFFF; assign b = 64'h345FFFFFFFFFFFFF;

    #10 $display("\n2**-836 * 2**-187:");
    #10 assign a = 64'h0BB0000000000000; assign b = 64'h3440000000000000;
    #10 assign a = 64'h0BBFFFFFFFFFFFFF; assign b = 64'h344FFFFFFFFFFFFF;

    #10 $display("\n2**-835 * 2**-188:");
    #10 assign a = 64'h0BC0000000000000; assign b = 64'h3430000000000000;
    #10 assign a = 64'h0BCFFFFFFFFFFFFF; assign b = 64'h343FFFFFFFFFFFFF;

    #10 $display("\n2**-834 * 2**-189:");
    #10 assign a = 64'h0BD0000000000000; assign b = 64'h3420000000000000;
    #10 assign a = 64'h0BDFFFFFFFFFFFFF; assign b = 64'h342FFFFFFFFFFFFF;

    #10 $display("\n2**-833 * 2**-190:");
    #10 assign a = 64'h0BE0000000000000; assign b = 64'h3410000000000000;
    #10 assign a = 64'h0BEFFFFFFFFFFFFF; assign b = 64'h341FFFFFFFFFFFFF;

    #10 $display("\n2**-832 * 2**-191:");
    #10 assign a = 64'h0BF0000000000000; assign b = 64'h3400000000000000;
    #10 assign a = 64'h0BFFFFFFFFFFFFFF; assign b = 64'h340FFFFFFFFFFFFF;

    #10 $display("\n2**-831 * 2**-192:");
    #10 assign a = 64'h0C00000000000000; assign b = 64'h33F0000000000000;
    #10 assign a = 64'h0C0FFFFFFFFFFFFF; assign b = 64'h33FFFFFFFFFFFFFF;

    #10 $display("\n2**-830 * 2**-193:");
    #10 assign a = 64'h0C10000000000000; assign b = 64'h33E0000000000000;
    #10 assign a = 64'h0C1FFFFFFFFFFFFF; assign b = 64'h33EFFFFFFFFFFFFF;

    #10 $display("\n2**-829 * 2**-194:");
    #10 assign a = 64'h0C20000000000000; assign b = 64'h33D0000000000000;
    #10 assign a = 64'h0C2FFFFFFFFFFFFF; assign b = 64'h33DFFFFFFFFFFFFF;

    #10 $display("\n2**-828 * 2**-195:");
    #10 assign a = 64'h0C30000000000000; assign b = 64'h33C0000000000000;
    #10 assign a = 64'h0C3FFFFFFFFFFFFF; assign b = 64'h33CFFFFFFFFFFFFF;

    #10 $display("\n2**-827 * 2**-196:");
    #10 assign a = 64'h0C40000000000000; assign b = 64'h33B0000000000000;
    #10 assign a = 64'h0C4FFFFFFFFFFFFF; assign b = 64'h33BFFFFFFFFFFFFF;

    #10 $display("\n2**-826 * 2**-197:");
    #10 assign a = 64'h0C50000000000000; assign b = 64'h33A0000000000000;
    #10 assign a = 64'h0C5FFFFFFFFFFFFF; assign b = 64'h33AFFFFFFFFFFFFF;

    #10 $display("\n2**-825 * 2**-198:");
    #10 assign a = 64'h0C60000000000000; assign b = 64'h3390000000000000;
    #10 assign a = 64'h0C6FFFFFFFFFFFFF; assign b = 64'h339FFFFFFFFFFFFF;

    #10 $display("\n2**-824 * 2**-199:");
    #10 assign a = 64'h0C70000000000000; assign b = 64'h3380000000000000;
    #10 assign a = 64'h0C7FFFFFFFFFFFFF; assign b = 64'h338FFFFFFFFFFFFF;

    #10 $display("\n2**-823 * 2**-200:");
    #10 assign a = 64'h0C80000000000000; assign b = 64'h3370000000000000;
    #10 assign a = 64'h0C8FFFFFFFFFFFFF; assign b = 64'h337FFFFFFFFFFFFF;

    #10 $display("\n2**-822 * 2**-201:");
    #10 assign a = 64'h0C90000000000000; assign b = 64'h3360000000000000;
    #10 assign a = 64'h0C9FFFFFFFFFFFFF; assign b = 64'h336FFFFFFFFFFFFF;

    #10 $display("\n2**-821 * 2**-202:");
    #10 assign a = 64'h0CA0000000000000; assign b = 64'h3350000000000000;
    #10 assign a = 64'h0CAFFFFFFFFFFFFF; assign b = 64'h335FFFFFFFFFFFFF;

    #10 $display("\n2**-820 * 2**-203:");
    #10 assign a = 64'h0CB0000000000000; assign b = 64'h3340000000000000;
    #10 assign a = 64'h0CBFFFFFFFFFFFFF; assign b = 64'h334FFFFFFFFFFFFF;

    #10 $display("\n2**-819 * 2**-204:");
    #10 assign a = 64'h0CC0000000000000; assign b = 64'h3330000000000000;
    #10 assign a = 64'h0CCFFFFFFFFFFFFF; assign b = 64'h333FFFFFFFFFFFFF;

    #10 $display("\n2**-818 * 2**-205:");
    #10 assign a = 64'h0CD0000000000000; assign b = 64'h3320000000000000;
    #10 assign a = 64'h0CDFFFFFFFFFFFFF; assign b = 64'h332FFFFFFFFFFFFF;

    #10 $display("\n2**-817 * 2**-206:");
    #10 assign a = 64'h0CE0000000000000; assign b = 64'h3310000000000000;
    #10 assign a = 64'h0CEFFFFFFFFFFFFF; assign b = 64'h331FFFFFFFFFFFFF;

    #10 $display("\n2**-816 * 2**-207:");
    #10 assign a = 64'h0CF0000000000000; assign b = 64'h3300000000000000;
    #10 assign a = 64'h0CFFFFFFFFFFFFFF; assign b = 64'h330FFFFFFFFFFFFF;

    #10 $display("\n2**-815 * 2**-208:");
    #10 assign a = 64'h0D00000000000000; assign b = 64'h32F0000000000000;
    #10 assign a = 64'h0D0FFFFFFFFFFFFF; assign b = 64'h32FFFFFFFFFFFFFF;

    #10 $display("\n2**-814 * 2**-209:");
    #10 assign a = 64'h0D10000000000000; assign b = 64'h32E0000000000000;
    #10 assign a = 64'h0D1FFFFFFFFFFFFF; assign b = 64'h32EFFFFFFFFFFFFF;

    #10 $display("\n2**-813 * 2**-210:");
    #10 assign a = 64'h0D20000000000000; assign b = 64'h32D0000000000000;
    #10 assign a = 64'h0D2FFFFFFFFFFFFF; assign b = 64'h32DFFFFFFFFFFFFF;

    #10 $display("\n2**-812 * 2**-211:");
    #10 assign a = 64'h0D30000000000000; assign b = 64'h32C0000000000000;
    #10 assign a = 64'h0D3FFFFFFFFFFFFF; assign b = 64'h32CFFFFFFFFFFFFF;

    #10 $display("\n2**-811 * 2**-212:");
    #10 assign a = 64'h0D40000000000000; assign b = 64'h32B0000000000000;
    #10 assign a = 64'h0D4FFFFFFFFFFFFF; assign b = 64'h32BFFFFFFFFFFFFF;

    #10 $display("\n2**-810 * 2**-213:");
    #10 assign a = 64'h0D50000000000000; assign b = 64'h32A0000000000000;
    #10 assign a = 64'h0D5FFFFFFFFFFFFF; assign b = 64'h32AFFFFFFFFFFFFF;

    #10 $display("\n2**-809 * 2**-214:");
    #10 assign a = 64'h0D60000000000000; assign b = 64'h3290000000000000;
    #10 assign a = 64'h0D6FFFFFFFFFFFFF; assign b = 64'h329FFFFFFFFFFFFF;

    #10 $display("\n2**-808 * 2**-215:");
    #10 assign a = 64'h0D70000000000000; assign b = 64'h3280000000000000;
    #10 assign a = 64'h0D7FFFFFFFFFFFFF; assign b = 64'h328FFFFFFFFFFFFF;

    #10 $display("\n2**-807 * 2**-216:");
    #10 assign a = 64'h0D80000000000000; assign b = 64'h3270000000000000;
    #10 assign a = 64'h0D8FFFFFFFFFFFFF; assign b = 64'h327FFFFFFFFFFFFF;

    #10 $display("\n2**-806 * 2**-217:");
    #10 assign a = 64'h0D90000000000000; assign b = 64'h3260000000000000;
    #10 assign a = 64'h0D9FFFFFFFFFFFFF; assign b = 64'h326FFFFFFFFFFFFF;

    #10 $display("\n2**-805 * 2**-218:");
    #10 assign a = 64'h0DA0000000000000; assign b = 64'h3250000000000000;
    #10 assign a = 64'h0DAFFFFFFFFFFFFF; assign b = 64'h325FFFFFFFFFFFFF;

    #10 $display("\n2**-804 * 2**-219:");
    #10 assign a = 64'h0DB0000000000000; assign b = 64'h3240000000000000;
    #10 assign a = 64'h0DBFFFFFFFFFFFFF; assign b = 64'h324FFFFFFFFFFFFF;

    #10 $display("\n2**-803 * 2**-220:");
    #10 assign a = 64'h0DC0000000000000; assign b = 64'h3230000000000000;
    #10 assign a = 64'h0DCFFFFFFFFFFFFF; assign b = 64'h323FFFFFFFFFFFFF;

    #10 $display("\n2**-802 * 2**-221:");
    #10 assign a = 64'h0DD0000000000000; assign b = 64'h3220000000000000;
    #10 assign a = 64'h0DDFFFFFFFFFFFFF; assign b = 64'h322FFFFFFFFFFFFF;

    #10 $display("\n2**-801 * 2**-222:");
    #10 assign a = 64'h0DE0000000000000; assign b = 64'h3210000000000000;
    #10 assign a = 64'h0DEFFFFFFFFFFFFF; assign b = 64'h321FFFFFFFFFFFFF;

    #10 $display("\n2**-800 * 2**-223:");
    #10 assign a = 64'h0DF0000000000000; assign b = 64'h3200000000000000;
    #10 assign a = 64'h0DFFFFFFFFFFFFFF; assign b = 64'h320FFFFFFFFFFFFF;

    #10 $display("\n2**-799 * 2**-224:");
    #10 assign a = 64'h0E00000000000000; assign b = 64'h31F0000000000000;
    #10 assign a = 64'h0E0FFFFFFFFFFFFF; assign b = 64'h31FFFFFFFFFFFFFF;

    #10 $display("\n2**-798 * 2**-225:");
    #10 assign a = 64'h0E10000000000000; assign b = 64'h31E0000000000000;
    #10 assign a = 64'h0E1FFFFFFFFFFFFF; assign b = 64'h31EFFFFFFFFFFFFF;

    #10 $display("\n2**-797 * 2**-226:");
    #10 assign a = 64'h0E20000000000000; assign b = 64'h31D0000000000000;
    #10 assign a = 64'h0E2FFFFFFFFFFFFF; assign b = 64'h31DFFFFFFFFFFFFF;

    #10 $display("\n2**-796 * 2**-227:");
    #10 assign a = 64'h0E30000000000000; assign b = 64'h31C0000000000000;
    #10 assign a = 64'h0E3FFFFFFFFFFFFF; assign b = 64'h31CFFFFFFFFFFFFF;

    #10 $display("\n2**-795 * 2**-228:");
    #10 assign a = 64'h0E40000000000000; assign b = 64'h31B0000000000000;
    #10 assign a = 64'h0E4FFFFFFFFFFFFF; assign b = 64'h31BFFFFFFFFFFFFF;

    #10 $display("\n2**-794 * 2**-229:");
    #10 assign a = 64'h0E50000000000000; assign b = 64'h31A0000000000000;
    #10 assign a = 64'h0E5FFFFFFFFFFFFF; assign b = 64'h31AFFFFFFFFFFFFF;

    #10 $display("\n2**-793 * 2**-230:");
    #10 assign a = 64'h0E60000000000000; assign b = 64'h3190000000000000;
    #10 assign a = 64'h0E6FFFFFFFFFFFFF; assign b = 64'h319FFFFFFFFFFFFF;

    #10 $display("\n2**-792 * 2**-231:");
    #10 assign a = 64'h0E70000000000000; assign b = 64'h3180000000000000;
    #10 assign a = 64'h0E7FFFFFFFFFFFFF; assign b = 64'h318FFFFFFFFFFFFF;

    #10 $display("\n2**-791 * 2**-232:");
    #10 assign a = 64'h0E80000000000000; assign b = 64'h3170000000000000;
    #10 assign a = 64'h0E8FFFFFFFFFFFFF; assign b = 64'h317FFFFFFFFFFFFF;

    #10 $display("\n2**-790 * 2**-233:");
    #10 assign a = 64'h0E90000000000000; assign b = 64'h3160000000000000;
    #10 assign a = 64'h0E9FFFFFFFFFFFFF; assign b = 64'h316FFFFFFFFFFFFF;

    #10 $display("\n2**-789 * 2**-234:");
    #10 assign a = 64'h0EA0000000000000; assign b = 64'h3150000000000000;
    #10 assign a = 64'h0EAFFFFFFFFFFFFF; assign b = 64'h315FFFFFFFFFFFFF;

    #10 $display("\n2**-788 * 2**-235:");
    #10 assign a = 64'h0EB0000000000000; assign b = 64'h3140000000000000;
    #10 assign a = 64'h0EBFFFFFFFFFFFFF; assign b = 64'h314FFFFFFFFFFFFF;

    #10 $display("\n2**-787 * 2**-236:");
    #10 assign a = 64'h0EC0000000000000; assign b = 64'h3130000000000000;
    #10 assign a = 64'h0ECFFFFFFFFFFFFF; assign b = 64'h313FFFFFFFFFFFFF;

    #10 $display("\n2**-786 * 2**-237:");
    #10 assign a = 64'h0ED0000000000000; assign b = 64'h3120000000000000;
    #10 assign a = 64'h0EDFFFFFFFFFFFFF; assign b = 64'h312FFFFFFFFFFFFF;

    #10 $display("\n2**-785 * 2**-238:");
    #10 assign a = 64'h0EE0000000000000; assign b = 64'h3110000000000000;
    #10 assign a = 64'h0EEFFFFFFFFFFFFF; assign b = 64'h311FFFFFFFFFFFFF;

    #10 $display("\n2**-784 * 2**-239:");
    #10 assign a = 64'h0EF0000000000000; assign b = 64'h3100000000000000;
    #10 assign a = 64'h0EFFFFFFFFFFFFFF; assign b = 64'h310FFFFFFFFFFFFF;

    #10 $display("\n2**-783 * 2**-240:");
    #10 assign a = 64'h0F00000000000000; assign b = 64'h30F0000000000000;
    #10 assign a = 64'h0F0FFFFFFFFFFFFF; assign b = 64'h30FFFFFFFFFFFFFF;

    #10 $display("\n2**-782 * 2**-241:");
    #10 assign a = 64'h0F10000000000000; assign b = 64'h30E0000000000000;
    #10 assign a = 64'h0F1FFFFFFFFFFFFF; assign b = 64'h30EFFFFFFFFFFFFF;

    #10 $display("\n2**-781 * 2**-242:");
    #10 assign a = 64'h0F20000000000000; assign b = 64'h30D0000000000000;
    #10 assign a = 64'h0F2FFFFFFFFFFFFF; assign b = 64'h30DFFFFFFFFFFFFF;

    #10 $display("\n2**-780 * 2**-243:");
    #10 assign a = 64'h0F30000000000000; assign b = 64'h30C0000000000000;
    #10 assign a = 64'h0F3FFFFFFFFFFFFF; assign b = 64'h30CFFFFFFFFFFFFF;

    #10 $display("\n2**-779 * 2**-244:");
    #10 assign a = 64'h0F40000000000000; assign b = 64'h30B0000000000000;
    #10 assign a = 64'h0F4FFFFFFFFFFFFF; assign b = 64'h30BFFFFFFFFFFFFF;

    #10 $display("\n2**-778 * 2**-245:");
    #10 assign a = 64'h0F50000000000000; assign b = 64'h30A0000000000000;
    #10 assign a = 64'h0F5FFFFFFFFFFFFF; assign b = 64'h30AFFFFFFFFFFFFF;

    #10 $display("\n2**-777 * 2**-246:");
    #10 assign a = 64'h0F60000000000000; assign b = 64'h3090000000000000;
    #10 assign a = 64'h0F6FFFFFFFFFFFFF; assign b = 64'h309FFFFFFFFFFFFF;

    #10 $display("\n2**-776 * 2**-247:");
    #10 assign a = 64'h0F70000000000000; assign b = 64'h3080000000000000;
    #10 assign a = 64'h0F7FFFFFFFFFFFFF; assign b = 64'h308FFFFFFFFFFFFF;

    #10 $display("\n2**-775 * 2**-248:");
    #10 assign a = 64'h0F80000000000000; assign b = 64'h3070000000000000;
    #10 assign a = 64'h0F8FFFFFFFFFFFFF; assign b = 64'h307FFFFFFFFFFFFF;

    #10 $display("\n2**-774 * 2**-249:");
    #10 assign a = 64'h0F90000000000000; assign b = 64'h3060000000000000;
    #10 assign a = 64'h0F9FFFFFFFFFFFFF; assign b = 64'h306FFFFFFFFFFFFF;

    #10 $display("\n2**-773 * 2**-250:");
    #10 assign a = 64'h0FA0000000000000; assign b = 64'h3050000000000000;
    #10 assign a = 64'h0FAFFFFFFFFFFFFF; assign b = 64'h305FFFFFFFFFFFFF;

    #10 $display("\n2**-772 * 2**-251:");
    #10 assign a = 64'h0FB0000000000000; assign b = 64'h3040000000000000;
    #10 assign a = 64'h0FBFFFFFFFFFFFFF; assign b = 64'h304FFFFFFFFFFFFF;

    #10 $display("\n2**-771 * 2**-252:");
    #10 assign a = 64'h0FC0000000000000; assign b = 64'h3030000000000000;
    #10 assign a = 64'h0FCFFFFFFFFFFFFF; assign b = 64'h303FFFFFFFFFFFFF;

    #10 $display("\n2**-770 * 2**-253:");
    #10 assign a = 64'h0FD0000000000000; assign b = 64'h3020000000000000;
    #10 assign a = 64'h0FDFFFFFFFFFFFFF; assign b = 64'h302FFFFFFFFFFFFF;

    #10 $display("\n2**-769 * 2**-254:");
    #10 assign a = 64'h0FE0000000000000; assign b = 64'h3010000000000000;
    #10 assign a = 64'h0FEFFFFFFFFFFFFF; assign b = 64'h301FFFFFFFFFFFFF;

    #10 $display("\n2**-768 * 2**-255:");
    #10 assign a = 64'h0FF0000000000000; assign b = 64'h3000000000000000;
    #10 assign a = 64'h0FFFFFFFFFFFFFFF; assign b = 64'h300FFFFFFFFFFFFF;

    #10 $display("\n2**-767 * 2**-256:");
    #10 assign a = 64'h1000000000000000; assign b = 64'h2FF0000000000000;
    #10 assign a = 64'h100FFFFFFFFFFFFF; assign b = 64'h2FFFFFFFFFFFFFFF;

    #10 $display("\n2**-766 * 2**-257:");
    #10 assign a = 64'h1010000000000000; assign b = 64'h2FE0000000000000;
    #10 assign a = 64'h101FFFFFFFFFFFFF; assign b = 64'h2FEFFFFFFFFFFFFF;

    #10 $display("\n2**-765 * 2**-258:");
    #10 assign a = 64'h1020000000000000; assign b = 64'h2FD0000000000000;
    #10 assign a = 64'h102FFFFFFFFFFFFF; assign b = 64'h2FDFFFFFFFFFFFFF;

    #10 $display("\n2**-764 * 2**-259:");
    #10 assign a = 64'h1030000000000000; assign b = 64'h2FC0000000000000;
    #10 assign a = 64'h103FFFFFFFFFFFFF; assign b = 64'h2FCFFFFFFFFFFFFF;

    #10 $display("\n2**-763 * 2**-260:");
    #10 assign a = 64'h1040000000000000; assign b = 64'h2FB0000000000000;
    #10 assign a = 64'h104FFFFFFFFFFFFF; assign b = 64'h2FBFFFFFFFFFFFFF;

    #10 $display("\n2**-762 * 2**-261:");
    #10 assign a = 64'h1050000000000000; assign b = 64'h2FA0000000000000;
    #10 assign a = 64'h105FFFFFFFFFFFFF; assign b = 64'h2FAFFFFFFFFFFFFF;

    #10 $display("\n2**-761 * 2**-262:");
    #10 assign a = 64'h1060000000000000; assign b = 64'h2F90000000000000;
    #10 assign a = 64'h106FFFFFFFFFFFFF; assign b = 64'h2F9FFFFFFFFFFFFF;

    #10 $display("\n2**-760 * 2**-263:");
    #10 assign a = 64'h1070000000000000; assign b = 64'h2F80000000000000;
    #10 assign a = 64'h107FFFFFFFFFFFFF; assign b = 64'h2F8FFFFFFFFFFFFF;

    #10 $display("\n2**-759 * 2**-264:");
    #10 assign a = 64'h1080000000000000; assign b = 64'h2F70000000000000;
    #10 assign a = 64'h108FFFFFFFFFFFFF; assign b = 64'h2F7FFFFFFFFFFFFF;

    #10 $display("\n2**-758 * 2**-265:");
    #10 assign a = 64'h1090000000000000; assign b = 64'h2F60000000000000;
    #10 assign a = 64'h109FFFFFFFFFFFFF; assign b = 64'h2F6FFFFFFFFFFFFF;

    #10 $display("\n2**-757 * 2**-266:");
    #10 assign a = 64'h10A0000000000000; assign b = 64'h2F50000000000000;
    #10 assign a = 64'h10AFFFFFFFFFFFFF; assign b = 64'h2F5FFFFFFFFFFFFF;

    #10 $display("\n2**-756 * 2**-267:");
    #10 assign a = 64'h10B0000000000000; assign b = 64'h2F40000000000000;
    #10 assign a = 64'h10BFFFFFFFFFFFFF; assign b = 64'h2F4FFFFFFFFFFFFF;

    #10 $display("\n2**-755 * 2**-268:");
    #10 assign a = 64'h10C0000000000000; assign b = 64'h2F30000000000000;
    #10 assign a = 64'h10CFFFFFFFFFFFFF; assign b = 64'h2F3FFFFFFFFFFFFF;

    #10 $display("\n2**-754 * 2**-269:");
    #10 assign a = 64'h10D0000000000000; assign b = 64'h2F20000000000000;
    #10 assign a = 64'h10DFFFFFFFFFFFFF; assign b = 64'h2F2FFFFFFFFFFFFF;

    #10 $display("\n2**-753 * 2**-270:");
    #10 assign a = 64'h10E0000000000000; assign b = 64'h2F10000000000000;
    #10 assign a = 64'h10EFFFFFFFFFFFFF; assign b = 64'h2F1FFFFFFFFFFFFF;

    #10 $display("\n2**-752 * 2**-271:");
    #10 assign a = 64'h10F0000000000000; assign b = 64'h2F00000000000000;
    #10 assign a = 64'h10FFFFFFFFFFFFFF; assign b = 64'h2F0FFFFFFFFFFFFF;

    #10 $display("\n2**-751 * 2**-272:");
    #10 assign a = 64'h1100000000000000; assign b = 64'h2EF0000000000000;
    #10 assign a = 64'h110FFFFFFFFFFFFF; assign b = 64'h2EFFFFFFFFFFFFFF;

    #10 $display("\n2**-750 * 2**-273:");
    #10 assign a = 64'h1110000000000000; assign b = 64'h2EE0000000000000;
    #10 assign a = 64'h111FFFFFFFFFFFFF; assign b = 64'h2EEFFFFFFFFFFFFF;

    #10 $display("\n2**-749 * 2**-274:");
    #10 assign a = 64'h1120000000000000; assign b = 64'h2ED0000000000000;
    #10 assign a = 64'h112FFFFFFFFFFFFF; assign b = 64'h2EDFFFFFFFFFFFFF;

    #10 $display("\n2**-748 * 2**-275:");
    #10 assign a = 64'h1130000000000000; assign b = 64'h2EC0000000000000;
    #10 assign a = 64'h113FFFFFFFFFFFFF; assign b = 64'h2ECFFFFFFFFFFFFF;

    #10 $display("\n2**-747 * 2**-276:");
    #10 assign a = 64'h1140000000000000; assign b = 64'h2EB0000000000000;
    #10 assign a = 64'h114FFFFFFFFFFFFF; assign b = 64'h2EBFFFFFFFFFFFFF;

    #10 $display("\n2**-746 * 2**-277:");
    #10 assign a = 64'h1150000000000000; assign b = 64'h2EA0000000000000;
    #10 assign a = 64'h115FFFFFFFFFFFFF; assign b = 64'h2EAFFFFFFFFFFFFF;

    #10 $display("\n2**-745 * 2**-278:");
    #10 assign a = 64'h1160000000000000; assign b = 64'h2E90000000000000;
    #10 assign a = 64'h116FFFFFFFFFFFFF; assign b = 64'h2E9FFFFFFFFFFFFF;

    #10 $display("\n2**-744 * 2**-279:");
    #10 assign a = 64'h1170000000000000; assign b = 64'h2E80000000000000;
    #10 assign a = 64'h117FFFFFFFFFFFFF; assign b = 64'h2E8FFFFFFFFFFFFF;

    #10 $display("\n2**-743 * 2**-280:");
    #10 assign a = 64'h1180000000000000; assign b = 64'h2E70000000000000;
    #10 assign a = 64'h118FFFFFFFFFFFFF; assign b = 64'h2E7FFFFFFFFFFFFF;

    #10 $display("\n2**-742 * 2**-281:");
    #10 assign a = 64'h1190000000000000; assign b = 64'h2E60000000000000;
    #10 assign a = 64'h119FFFFFFFFFFFFF; assign b = 64'h2E6FFFFFFFFFFFFF;

    #10 $display("\n2**-741 * 2**-282:");
    #10 assign a = 64'h11A0000000000000; assign b = 64'h2E50000000000000;
    #10 assign a = 64'h11AFFFFFFFFFFFFF; assign b = 64'h2E5FFFFFFFFFFFFF;

    #10 $display("\n2**-740 * 2**-283:");
    #10 assign a = 64'h11B0000000000000; assign b = 64'h2E40000000000000;
    #10 assign a = 64'h11BFFFFFFFFFFFFF; assign b = 64'h2E4FFFFFFFFFFFFF;

    #10 $display("\n2**-739 * 2**-284:");
    #10 assign a = 64'h11C0000000000000; assign b = 64'h2E30000000000000;
    #10 assign a = 64'h11CFFFFFFFFFFFFF; assign b = 64'h2E3FFFFFFFFFFFFF;

    #10 $display("\n2**-738 * 2**-285:");
    #10 assign a = 64'h11D0000000000000; assign b = 64'h2E20000000000000;
    #10 assign a = 64'h11DFFFFFFFFFFFFF; assign b = 64'h2E2FFFFFFFFFFFFF;

    #10 $display("\n2**-737 * 2**-286:");
    #10 assign a = 64'h11E0000000000000; assign b = 64'h2E10000000000000;
    #10 assign a = 64'h11EFFFFFFFFFFFFF; assign b = 64'h2E1FFFFFFFFFFFFF;

    #10 $display("\n2**-736 * 2**-287:");
    #10 assign a = 64'h11F0000000000000; assign b = 64'h2E00000000000000;
    #10 assign a = 64'h11FFFFFFFFFFFFFF; assign b = 64'h2E0FFFFFFFFFFFFF;

    #10 $display("\n2**-735 * 2**-288:");
    #10 assign a = 64'h1200000000000000; assign b = 64'h2DF0000000000000;
    #10 assign a = 64'h120FFFFFFFFFFFFF; assign b = 64'h2DFFFFFFFFFFFFFF;

    #10 $display("\n2**-734 * 2**-289:");
    #10 assign a = 64'h1210000000000000; assign b = 64'h2DE0000000000000;
    #10 assign a = 64'h121FFFFFFFFFFFFF; assign b = 64'h2DEFFFFFFFFFFFFF;

    #10 $display("\n2**-733 * 2**-290:");
    #10 assign a = 64'h1220000000000000; assign b = 64'h2DD0000000000000;
    #10 assign a = 64'h122FFFFFFFFFFFFF; assign b = 64'h2DDFFFFFFFFFFFFF;

    #10 $display("\n2**-732 * 2**-291:");
    #10 assign a = 64'h1230000000000000; assign b = 64'h2DC0000000000000;
    #10 assign a = 64'h123FFFFFFFFFFFFF; assign b = 64'h2DCFFFFFFFFFFFFF;

    #10 $display("\n2**-731 * 2**-292:");
    #10 assign a = 64'h1240000000000000; assign b = 64'h2DB0000000000000;
    #10 assign a = 64'h124FFFFFFFFFFFFF; assign b = 64'h2DBFFFFFFFFFFFFF;

    #10 $display("\n2**-730 * 2**-293:");
    #10 assign a = 64'h1250000000000000; assign b = 64'h2DA0000000000000;
    #10 assign a = 64'h125FFFFFFFFFFFFF; assign b = 64'h2DAFFFFFFFFFFFFF;

    #10 $display("\n2**-729 * 2**-294:");
    #10 assign a = 64'h1260000000000000; assign b = 64'h2D90000000000000;
    #10 assign a = 64'h126FFFFFFFFFFFFF; assign b = 64'h2D9FFFFFFFFFFFFF;

    #10 $display("\n2**-728 * 2**-295:");
    #10 assign a = 64'h1270000000000000; assign b = 64'h2D80000000000000;
    #10 assign a = 64'h127FFFFFFFFFFFFF; assign b = 64'h2D8FFFFFFFFFFFFF;

    #10 $display("\n2**-727 * 2**-296:");
    #10 assign a = 64'h1280000000000000; assign b = 64'h2D70000000000000;
    #10 assign a = 64'h128FFFFFFFFFFFFF; assign b = 64'h2D7FFFFFFFFFFFFF;

    #10 $display("\n2**-726 * 2**-297:");
    #10 assign a = 64'h1290000000000000; assign b = 64'h2D60000000000000;
    #10 assign a = 64'h129FFFFFFFFFFFFF; assign b = 64'h2D6FFFFFFFFFFFFF;

    #10 $display("\n2**-725 * 2**-298:");
    #10 assign a = 64'h12A0000000000000; assign b = 64'h2D50000000000000;
    #10 assign a = 64'h12AFFFFFFFFFFFFF; assign b = 64'h2D5FFFFFFFFFFFFF;

    #10 $display("\n2**-724 * 2**-299:");
    #10 assign a = 64'h12B0000000000000; assign b = 64'h2D40000000000000;
    #10 assign a = 64'h12BFFFFFFFFFFFFF; assign b = 64'h2D4FFFFFFFFFFFFF;

    #10 $display("\n2**-723 * 2**-300:");
    #10 assign a = 64'h12C0000000000000; assign b = 64'h2D30000000000000;
    #10 assign a = 64'h12CFFFFFFFFFFFFF; assign b = 64'h2D3FFFFFFFFFFFFF;

    #10 $display("\n2**-722 * 2**-301:");
    #10 assign a = 64'h12D0000000000000; assign b = 64'h2D20000000000000;
    #10 assign a = 64'h12DFFFFFFFFFFFFF; assign b = 64'h2D2FFFFFFFFFFFFF;

    #10 $display("\n2**-721 * 2**-302:");
    #10 assign a = 64'h12E0000000000000; assign b = 64'h2D10000000000000;
    #10 assign a = 64'h12EFFFFFFFFFFFFF; assign b = 64'h2D1FFFFFFFFFFFFF;

    #10 $display("\n2**-720 * 2**-303:");
    #10 assign a = 64'h12F0000000000000; assign b = 64'h2D00000000000000;
    #10 assign a = 64'h12FFFFFFFFFFFFFF; assign b = 64'h2D0FFFFFFFFFFFFF;

    #10 $display("\n2**-719 * 2**-304:");
    #10 assign a = 64'h1300000000000000; assign b = 64'h2CF0000000000000;
    #10 assign a = 64'h130FFFFFFFFFFFFF; assign b = 64'h2CFFFFFFFFFFFFFF;

    #10 $display("\n2**-718 * 2**-305:");
    #10 assign a = 64'h1310000000000000; assign b = 64'h2CE0000000000000;
    #10 assign a = 64'h131FFFFFFFFFFFFF; assign b = 64'h2CEFFFFFFFFFFFFF;

    #10 $display("\n2**-717 * 2**-306:");
    #10 assign a = 64'h1320000000000000; assign b = 64'h2CD0000000000000;
    #10 assign a = 64'h132FFFFFFFFFFFFF; assign b = 64'h2CDFFFFFFFFFFFFF;

    #10 $display("\n2**-716 * 2**-307:");
    #10 assign a = 64'h1330000000000000; assign b = 64'h2CC0000000000000;
    #10 assign a = 64'h133FFFFFFFFFFFFF; assign b = 64'h2CCFFFFFFFFFFFFF;

    #10 $display("\n2**-715 * 2**-308:");
    #10 assign a = 64'h1340000000000000; assign b = 64'h2CB0000000000000;
    #10 assign a = 64'h134FFFFFFFFFFFFF; assign b = 64'h2CBFFFFFFFFFFFFF;

    #10 $display("\n2**-714 * 2**-309:");
    #10 assign a = 64'h1350000000000000; assign b = 64'h2CA0000000000000;
    #10 assign a = 64'h135FFFFFFFFFFFFF; assign b = 64'h2CAFFFFFFFFFFFFF;

    #10 $display("\n2**-713 * 2**-310:");
    #10 assign a = 64'h1360000000000000; assign b = 64'h2C90000000000000;
    #10 assign a = 64'h136FFFFFFFFFFFFF; assign b = 64'h2C9FFFFFFFFFFFFF;

    #10 $display("\n2**-712 * 2**-311:");
    #10 assign a = 64'h1370000000000000; assign b = 64'h2C80000000000000;
    #10 assign a = 64'h137FFFFFFFFFFFFF; assign b = 64'h2C8FFFFFFFFFFFFF;

    #10 $display("\n2**-711 * 2**-312:");
    #10 assign a = 64'h1380000000000000; assign b = 64'h2C70000000000000;
    #10 assign a = 64'h138FFFFFFFFFFFFF; assign b = 64'h2C7FFFFFFFFFFFFF;

    #10 $display("\n2**-710 * 2**-313:");
    #10 assign a = 64'h1390000000000000; assign b = 64'h2C60000000000000;
    #10 assign a = 64'h139FFFFFFFFFFFFF; assign b = 64'h2C6FFFFFFFFFFFFF;

    #10 $display("\n2**-709 * 2**-314:");
    #10 assign a = 64'h13A0000000000000; assign b = 64'h2C50000000000000;
    #10 assign a = 64'h13AFFFFFFFFFFFFF; assign b = 64'h2C5FFFFFFFFFFFFF;

    #10 $display("\n2**-708 * 2**-315:");
    #10 assign a = 64'h13B0000000000000; assign b = 64'h2C40000000000000;
    #10 assign a = 64'h13BFFFFFFFFFFFFF; assign b = 64'h2C4FFFFFFFFFFFFF;

    #10 $display("\n2**-707 * 2**-316:");
    #10 assign a = 64'h13C0000000000000; assign b = 64'h2C30000000000000;
    #10 assign a = 64'h13CFFFFFFFFFFFFF; assign b = 64'h2C3FFFFFFFFFFFFF;

    #10 $display("\n2**-706 * 2**-317:");
    #10 assign a = 64'h13D0000000000000; assign b = 64'h2C20000000000000;
    #10 assign a = 64'h13DFFFFFFFFFFFFF; assign b = 64'h2C2FFFFFFFFFFFFF;

    #10 $display("\n2**-705 * 2**-318:");
    #10 assign a = 64'h13E0000000000000; assign b = 64'h2C10000000000000;
    #10 assign a = 64'h13EFFFFFFFFFFFFF; assign b = 64'h2C1FFFFFFFFFFFFF;

    #10 $display("\n2**-704 * 2**-319:");
    #10 assign a = 64'h13F0000000000000; assign b = 64'h2C00000000000000;
    #10 assign a = 64'h13FFFFFFFFFFFFFF; assign b = 64'h2C0FFFFFFFFFFFFF;

    #10 $display("\n2**-703 * 2**-320:");
    #10 assign a = 64'h1400000000000000; assign b = 64'h2BF0000000000000;
    #10 assign a = 64'h140FFFFFFFFFFFFF; assign b = 64'h2BFFFFFFFFFFFFFF;

    #10 $display("\n2**-702 * 2**-321:");
    #10 assign a = 64'h1410000000000000; assign b = 64'h2BE0000000000000;
    #10 assign a = 64'h141FFFFFFFFFFFFF; assign b = 64'h2BEFFFFFFFFFFFFF;

    #10 $display("\n2**-701 * 2**-322:");
    #10 assign a = 64'h1420000000000000; assign b = 64'h2BD0000000000000;
    #10 assign a = 64'h142FFFFFFFFFFFFF; assign b = 64'h2BDFFFFFFFFFFFFF;

    #10 $display("\n2**-700 * 2**-323:");
    #10 assign a = 64'h1430000000000000; assign b = 64'h2BC0000000000000;
    #10 assign a = 64'h143FFFFFFFFFFFFF; assign b = 64'h2BCFFFFFFFFFFFFF;

    #10 $display("\n2**-699 * 2**-324:");
    #10 assign a = 64'h1440000000000000; assign b = 64'h2BB0000000000000;
    #10 assign a = 64'h144FFFFFFFFFFFFF; assign b = 64'h2BBFFFFFFFFFFFFF;

    #10 $display("\n2**-698 * 2**-325:");
    #10 assign a = 64'h1450000000000000; assign b = 64'h2BA0000000000000;
    #10 assign a = 64'h145FFFFFFFFFFFFF; assign b = 64'h2BAFFFFFFFFFFFFF;

    #10 $display("\n2**-697 * 2**-326:");
    #10 assign a = 64'h1460000000000000; assign b = 64'h2B90000000000000;
    #10 assign a = 64'h146FFFFFFFFFFFFF; assign b = 64'h2B9FFFFFFFFFFFFF;

    #10 $display("\n2**-696 * 2**-327:");
    #10 assign a = 64'h1470000000000000; assign b = 64'h2B80000000000000;
    #10 assign a = 64'h147FFFFFFFFFFFFF; assign b = 64'h2B8FFFFFFFFFFFFF;

    #10 $display("\n2**-695 * 2**-328:");
    #10 assign a = 64'h1480000000000000; assign b = 64'h2B70000000000000;
    #10 assign a = 64'h148FFFFFFFFFFFFF; assign b = 64'h2B7FFFFFFFFFFFFF;

    #10 $display("\n2**-694 * 2**-329:");
    #10 assign a = 64'h1490000000000000; assign b = 64'h2B60000000000000;
    #10 assign a = 64'h149FFFFFFFFFFFFF; assign b = 64'h2B6FFFFFFFFFFFFF;

    #10 $display("\n2**-693 * 2**-330:");
    #10 assign a = 64'h14A0000000000000; assign b = 64'h2B50000000000000;
    #10 assign a = 64'h14AFFFFFFFFFFFFF; assign b = 64'h2B5FFFFFFFFFFFFF;

    #10 $display("\n2**-692 * 2**-331:");
    #10 assign a = 64'h14B0000000000000; assign b = 64'h2B40000000000000;
    #10 assign a = 64'h14BFFFFFFFFFFFFF; assign b = 64'h2B4FFFFFFFFFFFFF;

    #10 $display("\n2**-691 * 2**-332:");
    #10 assign a = 64'h14C0000000000000; assign b = 64'h2B30000000000000;
    #10 assign a = 64'h14CFFFFFFFFFFFFF; assign b = 64'h2B3FFFFFFFFFFFFF;

    #10 $display("\n2**-690 * 2**-333:");
    #10 assign a = 64'h14D0000000000000; assign b = 64'h2B20000000000000;
    #10 assign a = 64'h14DFFFFFFFFFFFFF; assign b = 64'h2B2FFFFFFFFFFFFF;

    #10 $display("\n2**-689 * 2**-334:");
    #10 assign a = 64'h14E0000000000000; assign b = 64'h2B10000000000000;
    #10 assign a = 64'h14EFFFFFFFFFFFFF; assign b = 64'h2B1FFFFFFFFFFFFF;

    #10 $display("\n2**-688 * 2**-335:");
    #10 assign a = 64'h14F0000000000000; assign b = 64'h2B00000000000000;
    #10 assign a = 64'h14FFFFFFFFFFFFFF; assign b = 64'h2B0FFFFFFFFFFFFF;

    #10 $display("\n2**-687 * 2**-336:");
    #10 assign a = 64'h1500000000000000; assign b = 64'h2AF0000000000000;
    #10 assign a = 64'h150FFFFFFFFFFFFF; assign b = 64'h2AFFFFFFFFFFFFFF;

    #10 $display("\n2**-686 * 2**-337:");
    #10 assign a = 64'h1510000000000000; assign b = 64'h2AE0000000000000;
    #10 assign a = 64'h151FFFFFFFFFFFFF; assign b = 64'h2AEFFFFFFFFFFFFF;

    #10 $display("\n2**-685 * 2**-338:");
    #10 assign a = 64'h1520000000000000; assign b = 64'h2AD0000000000000;
    #10 assign a = 64'h152FFFFFFFFFFFFF; assign b = 64'h2ADFFFFFFFFFFFFF;

    #10 $display("\n2**-684 * 2**-339:");
    #10 assign a = 64'h1530000000000000; assign b = 64'h2AC0000000000000;
    #10 assign a = 64'h153FFFFFFFFFFFFF; assign b = 64'h2ACFFFFFFFFFFFFF;

    #10 $display("\n2**-683 * 2**-340:");
    #10 assign a = 64'h1540000000000000; assign b = 64'h2AB0000000000000;
    #10 assign a = 64'h154FFFFFFFFFFFFF; assign b = 64'h2ABFFFFFFFFFFFFF;

    #10 $display("\n2**-682 * 2**-341:");
    #10 assign a = 64'h1550000000000000; assign b = 64'h2AA0000000000000;
    #10 assign a = 64'h155FFFFFFFFFFFFF; assign b = 64'h2AAFFFFFFFFFFFFF;

    #10 $display("\n2**-681 * 2**-342:");
    #10 assign a = 64'h1560000000000000; assign b = 64'h2A90000000000000;
    #10 assign a = 64'h156FFFFFFFFFFFFF; assign b = 64'h2A9FFFFFFFFFFFFF;

    #10 $display("\n2**-680 * 2**-343:");
    #10 assign a = 64'h1570000000000000; assign b = 64'h2A80000000000000;
    #10 assign a = 64'h157FFFFFFFFFFFFF; assign b = 64'h2A8FFFFFFFFFFFFF;

    #10 $display("\n2**-679 * 2**-344:");
    #10 assign a = 64'h1580000000000000; assign b = 64'h2A70000000000000;
    #10 assign a = 64'h158FFFFFFFFFFFFF; assign b = 64'h2A7FFFFFFFFFFFFF;

    #10 $display("\n2**-678 * 2**-345:");
    #10 assign a = 64'h1590000000000000; assign b = 64'h2A60000000000000;
    #10 assign a = 64'h159FFFFFFFFFFFFF; assign b = 64'h2A6FFFFFFFFFFFFF;

    #10 $display("\n2**-677 * 2**-346:");
    #10 assign a = 64'h15A0000000000000; assign b = 64'h2A50000000000000;
    #10 assign a = 64'h15AFFFFFFFFFFFFF; assign b = 64'h2A5FFFFFFFFFFFFF;

    #10 $display("\n2**-676 * 2**-347:");
    #10 assign a = 64'h15B0000000000000; assign b = 64'h2A40000000000000;
    #10 assign a = 64'h15BFFFFFFFFFFFFF; assign b = 64'h2A4FFFFFFFFFFFFF;

    #10 $display("\n2**-675 * 2**-348:");
    #10 assign a = 64'h15C0000000000000; assign b = 64'h2A30000000000000;
    #10 assign a = 64'h15CFFFFFFFFFFFFF; assign b = 64'h2A3FFFFFFFFFFFFF;

    #10 $display("\n2**-674 * 2**-349:");
    #10 assign a = 64'h15D0000000000000; assign b = 64'h2A20000000000000;
    #10 assign a = 64'h15DFFFFFFFFFFFFF; assign b = 64'h2A2FFFFFFFFFFFFF;

    #10 $display("\n2**-673 * 2**-350:");
    #10 assign a = 64'h15E0000000000000; assign b = 64'h2A10000000000000;
    #10 assign a = 64'h15EFFFFFFFFFFFFF; assign b = 64'h2A1FFFFFFFFFFFFF;

    #10 $display("\n2**-672 * 2**-351:");
    #10 assign a = 64'h15F0000000000000; assign b = 64'h2A00000000000000;
    #10 assign a = 64'h15FFFFFFFFFFFFFF; assign b = 64'h2A0FFFFFFFFFFFFF;

    #10 $display("\n2**-671 * 2**-352:");
    #10 assign a = 64'h1600000000000000; assign b = 64'h29F0000000000000;
    #10 assign a = 64'h160FFFFFFFFFFFFF; assign b = 64'h29FFFFFFFFFFFFFF;

    #10 $display("\n2**-670 * 2**-353:");
    #10 assign a = 64'h1610000000000000; assign b = 64'h29E0000000000000;
    #10 assign a = 64'h161FFFFFFFFFFFFF; assign b = 64'h29EFFFFFFFFFFFFF;

    #10 $display("\n2**-669 * 2**-354:");
    #10 assign a = 64'h1620000000000000; assign b = 64'h29D0000000000000;
    #10 assign a = 64'h162FFFFFFFFFFFFF; assign b = 64'h29DFFFFFFFFFFFFF;

    #10 $display("\n2**-668 * 2**-355:");
    #10 assign a = 64'h1630000000000000; assign b = 64'h29C0000000000000;
    #10 assign a = 64'h163FFFFFFFFFFFFF; assign b = 64'h29CFFFFFFFFFFFFF;

    #10 $display("\n2**-667 * 2**-356:");
    #10 assign a = 64'h1640000000000000; assign b = 64'h29B0000000000000;
    #10 assign a = 64'h164FFFFFFFFFFFFF; assign b = 64'h29BFFFFFFFFFFFFF;

    #10 $display("\n2**-666 * 2**-357:");
    #10 assign a = 64'h1650000000000000; assign b = 64'h29A0000000000000;
    #10 assign a = 64'h165FFFFFFFFFFFFF; assign b = 64'h29AFFFFFFFFFFFFF;

    #10 $display("\n2**-665 * 2**-358:");
    #10 assign a = 64'h1660000000000000; assign b = 64'h2990000000000000;
    #10 assign a = 64'h166FFFFFFFFFFFFF; assign b = 64'h299FFFFFFFFFFFFF;

    #10 $display("\n2**-664 * 2**-359:");
    #10 assign a = 64'h1670000000000000; assign b = 64'h2980000000000000;
    #10 assign a = 64'h167FFFFFFFFFFFFF; assign b = 64'h298FFFFFFFFFFFFF;

    #10 $display("\n2**-663 * 2**-360:");
    #10 assign a = 64'h1680000000000000; assign b = 64'h2970000000000000;
    #10 assign a = 64'h168FFFFFFFFFFFFF; assign b = 64'h297FFFFFFFFFFFFF;

    #10 $display("\n2**-662 * 2**-361:");
    #10 assign a = 64'h1690000000000000; assign b = 64'h2960000000000000;
    #10 assign a = 64'h169FFFFFFFFFFFFF; assign b = 64'h296FFFFFFFFFFFFF;

    #10 $display("\n2**-661 * 2**-362:");
    #10 assign a = 64'h16A0000000000000; assign b = 64'h2950000000000000;
    #10 assign a = 64'h16AFFFFFFFFFFFFF; assign b = 64'h295FFFFFFFFFFFFF;

    #10 $display("\n2**-660 * 2**-363:");
    #10 assign a = 64'h16B0000000000000; assign b = 64'h2940000000000000;
    #10 assign a = 64'h16BFFFFFFFFFFFFF; assign b = 64'h294FFFFFFFFFFFFF;

    #10 $display("\n2**-659 * 2**-364:");
    #10 assign a = 64'h16C0000000000000; assign b = 64'h2930000000000000;
    #10 assign a = 64'h16CFFFFFFFFFFFFF; assign b = 64'h293FFFFFFFFFFFFF;

    #10 $display("\n2**-658 * 2**-365:");
    #10 assign a = 64'h16D0000000000000; assign b = 64'h2920000000000000;
    #10 assign a = 64'h16DFFFFFFFFFFFFF; assign b = 64'h292FFFFFFFFFFFFF;

    #10 $display("\n2**-657 * 2**-366:");
    #10 assign a = 64'h16E0000000000000; assign b = 64'h2910000000000000;
    #10 assign a = 64'h16EFFFFFFFFFFFFF; assign b = 64'h291FFFFFFFFFFFFF;

    #10 $display("\n2**-656 * 2**-367:");
    #10 assign a = 64'h16F0000000000000; assign b = 64'h2900000000000000;
    #10 assign a = 64'h16FFFFFFFFFFFFFF; assign b = 64'h290FFFFFFFFFFFFF;

    #10 $display("\n2**-655 * 2**-368:");
    #10 assign a = 64'h1700000000000000; assign b = 64'h28F0000000000000;
    #10 assign a = 64'h170FFFFFFFFFFFFF; assign b = 64'h28FFFFFFFFFFFFFF;

    #10 $display("\n2**-654 * 2**-369:");
    #10 assign a = 64'h1710000000000000; assign b = 64'h28E0000000000000;
    #10 assign a = 64'h171FFFFFFFFFFFFF; assign b = 64'h28EFFFFFFFFFFFFF;

    #10 $display("\n2**-653 * 2**-370:");
    #10 assign a = 64'h1720000000000000; assign b = 64'h28D0000000000000;
    #10 assign a = 64'h172FFFFFFFFFFFFF; assign b = 64'h28DFFFFFFFFFFFFF;

    #10 $display("\n2**-652 * 2**-371:");
    #10 assign a = 64'h1730000000000000; assign b = 64'h28C0000000000000;
    #10 assign a = 64'h173FFFFFFFFFFFFF; assign b = 64'h28CFFFFFFFFFFFFF;

    #10 $display("\n2**-651 * 2**-372:");
    #10 assign a = 64'h1740000000000000; assign b = 64'h28B0000000000000;
    #10 assign a = 64'h174FFFFFFFFFFFFF; assign b = 64'h28BFFFFFFFFFFFFF;

    #10 $display("\n2**-650 * 2**-373:");
    #10 assign a = 64'h1750000000000000; assign b = 64'h28A0000000000000;
    #10 assign a = 64'h175FFFFFFFFFFFFF; assign b = 64'h28AFFFFFFFFFFFFF;

    #10 $display("\n2**-649 * 2**-374:");
    #10 assign a = 64'h1760000000000000; assign b = 64'h2890000000000000;
    #10 assign a = 64'h176FFFFFFFFFFFFF; assign b = 64'h289FFFFFFFFFFFFF;

    #10 $display("\n2**-648 * 2**-375:");
    #10 assign a = 64'h1770000000000000; assign b = 64'h2880000000000000;
    #10 assign a = 64'h177FFFFFFFFFFFFF; assign b = 64'h288FFFFFFFFFFFFF;

    #10 $display("\n2**-647 * 2**-376:");
    #10 assign a = 64'h1780000000000000; assign b = 64'h2870000000000000;
    #10 assign a = 64'h178FFFFFFFFFFFFF; assign b = 64'h287FFFFFFFFFFFFF;

    #10 $display("\n2**-646 * 2**-377:");
    #10 assign a = 64'h1790000000000000; assign b = 64'h2860000000000000;
    #10 assign a = 64'h179FFFFFFFFFFFFF; assign b = 64'h286FFFFFFFFFFFFF;

    #10 $display("\n2**-645 * 2**-378:");
    #10 assign a = 64'h17A0000000000000; assign b = 64'h2850000000000000;
    #10 assign a = 64'h17AFFFFFFFFFFFFF; assign b = 64'h285FFFFFFFFFFFFF;

    #10 $display("\n2**-644 * 2**-379:");
    #10 assign a = 64'h17B0000000000000; assign b = 64'h2840000000000000;
    #10 assign a = 64'h17BFFFFFFFFFFFFF; assign b = 64'h284FFFFFFFFFFFFF;

    #10 $display("\n2**-643 * 2**-380:");
    #10 assign a = 64'h17C0000000000000; assign b = 64'h2830000000000000;
    #10 assign a = 64'h17CFFFFFFFFFFFFF; assign b = 64'h283FFFFFFFFFFFFF;

    #10 $display("\n2**-642 * 2**-381:");
    #10 assign a = 64'h17D0000000000000; assign b = 64'h2820000000000000;
    #10 assign a = 64'h17DFFFFFFFFFFFFF; assign b = 64'h282FFFFFFFFFFFFF;

    #10 $display("\n2**-641 * 2**-382:");
    #10 assign a = 64'h17E0000000000000; assign b = 64'h2810000000000000;
    #10 assign a = 64'h17EFFFFFFFFFFFFF; assign b = 64'h281FFFFFFFFFFFFF;

    #10 $display("\n2**-640 * 2**-383:");
    #10 assign a = 64'h17F0000000000000; assign b = 64'h2800000000000000;
    #10 assign a = 64'h17FFFFFFFFFFFFFF; assign b = 64'h280FFFFFFFFFFFFF;

    #10 $display("\n2**-639 * 2**-384:");
    #10 assign a = 64'h1800000000000000; assign b = 64'h27F0000000000000;
    #10 assign a = 64'h180FFFFFFFFFFFFF; assign b = 64'h27FFFFFFFFFFFFFF;

    #10 $display("\n2**-638 * 2**-385:");
    #10 assign a = 64'h1810000000000000; assign b = 64'h27E0000000000000;
    #10 assign a = 64'h181FFFFFFFFFFFFF; assign b = 64'h27EFFFFFFFFFFFFF;

    #10 $display("\n2**-637 * 2**-386:");
    #10 assign a = 64'h1820000000000000; assign b = 64'h27D0000000000000;
    #10 assign a = 64'h182FFFFFFFFFFFFF; assign b = 64'h27DFFFFFFFFFFFFF;

    #10 $display("\n2**-636 * 2**-387:");
    #10 assign a = 64'h1830000000000000; assign b = 64'h27C0000000000000;
    #10 assign a = 64'h183FFFFFFFFFFFFF; assign b = 64'h27CFFFFFFFFFFFFF;

    #10 $display("\n2**-635 * 2**-388:");
    #10 assign a = 64'h1840000000000000; assign b = 64'h27B0000000000000;
    #10 assign a = 64'h184FFFFFFFFFFFFF; assign b = 64'h27BFFFFFFFFFFFFF;

    #10 $display("\n2**-634 * 2**-389:");
    #10 assign a = 64'h1850000000000000; assign b = 64'h27A0000000000000;
    #10 assign a = 64'h185FFFFFFFFFFFFF; assign b = 64'h27AFFFFFFFFFFFFF;

    #10 $display("\n2**-633 * 2**-390:");
    #10 assign a = 64'h1860000000000000; assign b = 64'h2790000000000000;
    #10 assign a = 64'h186FFFFFFFFFFFFF; assign b = 64'h279FFFFFFFFFFFFF;

    #10 $display("\n2**-632 * 2**-391:");
    #10 assign a = 64'h1870000000000000; assign b = 64'h2780000000000000;
    #10 assign a = 64'h187FFFFFFFFFFFFF; assign b = 64'h278FFFFFFFFFFFFF;

    #10 $display("\n2**-631 * 2**-392:");
    #10 assign a = 64'h1880000000000000; assign b = 64'h2770000000000000;
    #10 assign a = 64'h188FFFFFFFFFFFFF; assign b = 64'h277FFFFFFFFFFFFF;

    #10 $display("\n2**-630 * 2**-393:");
    #10 assign a = 64'h1890000000000000; assign b = 64'h2760000000000000;
    #10 assign a = 64'h189FFFFFFFFFFFFF; assign b = 64'h276FFFFFFFFFFFFF;

    #10 $display("\n2**-629 * 2**-394:");
    #10 assign a = 64'h18A0000000000000; assign b = 64'h2750000000000000;
    #10 assign a = 64'h18AFFFFFFFFFFFFF; assign b = 64'h275FFFFFFFFFFFFF;

    #10 $display("\n2**-628 * 2**-395:");
    #10 assign a = 64'h18B0000000000000; assign b = 64'h2740000000000000;
    #10 assign a = 64'h18BFFFFFFFFFFFFF; assign b = 64'h274FFFFFFFFFFFFF;

    #10 $display("\n2**-627 * 2**-396:");
    #10 assign a = 64'h18C0000000000000; assign b = 64'h2730000000000000;
    #10 assign a = 64'h18CFFFFFFFFFFFFF; assign b = 64'h273FFFFFFFFFFFFF;

    #10 $display("\n2**-626 * 2**-397:");
    #10 assign a = 64'h18D0000000000000; assign b = 64'h2720000000000000;
    #10 assign a = 64'h18DFFFFFFFFFFFFF; assign b = 64'h272FFFFFFFFFFFFF;

    #10 $display("\n2**-625 * 2**-398:");
    #10 assign a = 64'h18E0000000000000; assign b = 64'h2710000000000000;
    #10 assign a = 64'h18EFFFFFFFFFFFFF; assign b = 64'h271FFFFFFFFFFFFF;

    #10 $display("\n2**-624 * 2**-399:");
    #10 assign a = 64'h18F0000000000000; assign b = 64'h2700000000000000;
    #10 assign a = 64'h18FFFFFFFFFFFFFF; assign b = 64'h270FFFFFFFFFFFFF;

    #10 $display("\n2**-623 * 2**-400:");
    #10 assign a = 64'h1900000000000000; assign b = 64'h26F0000000000000;
    #10 assign a = 64'h190FFFFFFFFFFFFF; assign b = 64'h26FFFFFFFFFFFFFF;

    #10 $display("\n2**-622 * 2**-401:");
    #10 assign a = 64'h1910000000000000; assign b = 64'h26E0000000000000;
    #10 assign a = 64'h191FFFFFFFFFFFFF; assign b = 64'h26EFFFFFFFFFFFFF;

    #10 $display("\n2**-621 * 2**-402:");
    #10 assign a = 64'h1920000000000000; assign b = 64'h26D0000000000000;
    #10 assign a = 64'h192FFFFFFFFFFFFF; assign b = 64'h26DFFFFFFFFFFFFF;

    #10 $display("\n2**-620 * 2**-403:");
    #10 assign a = 64'h1930000000000000; assign b = 64'h26C0000000000000;
    #10 assign a = 64'h193FFFFFFFFFFFFF; assign b = 64'h26CFFFFFFFFFFFFF;

    #10 $display("\n2**-619 * 2**-404:");
    #10 assign a = 64'h1940000000000000; assign b = 64'h26B0000000000000;
    #10 assign a = 64'h194FFFFFFFFFFFFF; assign b = 64'h26BFFFFFFFFFFFFF;

    #10 $display("\n2**-618 * 2**-405:");
    #10 assign a = 64'h1950000000000000; assign b = 64'h26A0000000000000;
    #10 assign a = 64'h195FFFFFFFFFFFFF; assign b = 64'h26AFFFFFFFFFFFFF;

    #10 $display("\n2**-617 * 2**-406:");
    #10 assign a = 64'h1960000000000000; assign b = 64'h2690000000000000;
    #10 assign a = 64'h196FFFFFFFFFFFFF; assign b = 64'h269FFFFFFFFFFFFF;

    #10 $display("\n2**-616 * 2**-407:");
    #10 assign a = 64'h1970000000000000; assign b = 64'h2680000000000000;
    #10 assign a = 64'h197FFFFFFFFFFFFF; assign b = 64'h268FFFFFFFFFFFFF;

    #10 $display("\n2**-615 * 2**-408:");
    #10 assign a = 64'h1980000000000000; assign b = 64'h2670000000000000;
    #10 assign a = 64'h198FFFFFFFFFFFFF; assign b = 64'h267FFFFFFFFFFFFF;

    #10 $display("\n2**-614 * 2**-409:");
    #10 assign a = 64'h1990000000000000; assign b = 64'h2660000000000000;
    #10 assign a = 64'h199FFFFFFFFFFFFF; assign b = 64'h266FFFFFFFFFFFFF;

    #10 $display("\n2**-613 * 2**-410:");
    #10 assign a = 64'h19A0000000000000; assign b = 64'h2650000000000000;
    #10 assign a = 64'h19AFFFFFFFFFFFFF; assign b = 64'h265FFFFFFFFFFFFF;

    #10 $display("\n2**-612 * 2**-411:");
    #10 assign a = 64'h19B0000000000000; assign b = 64'h2640000000000000;
    #10 assign a = 64'h19BFFFFFFFFFFFFF; assign b = 64'h264FFFFFFFFFFFFF;

    #10 $display("\n2**-611 * 2**-412:");
    #10 assign a = 64'h19C0000000000000; assign b = 64'h2630000000000000;
    #10 assign a = 64'h19CFFFFFFFFFFFFF; assign b = 64'h263FFFFFFFFFFFFF;

    #10 $display("\n2**-610 * 2**-413:");
    #10 assign a = 64'h19D0000000000000; assign b = 64'h2620000000000000;
    #10 assign a = 64'h19DFFFFFFFFFFFFF; assign b = 64'h262FFFFFFFFFFFFF;

    #10 $display("\n2**-609 * 2**-414:");
    #10 assign a = 64'h19E0000000000000; assign b = 64'h2610000000000000;
    #10 assign a = 64'h19EFFFFFFFFFFFFF; assign b = 64'h261FFFFFFFFFFFFF;

    #10 $display("\n2**-608 * 2**-415:");
    #10 assign a = 64'h19F0000000000000; assign b = 64'h2600000000000000;
    #10 assign a = 64'h19FFFFFFFFFFFFFF; assign b = 64'h260FFFFFFFFFFFFF;

    #10 $display("\n2**-607 * 2**-416:");
    #10 assign a = 64'h1A00000000000000; assign b = 64'h25F0000000000000;
    #10 assign a = 64'h1A0FFFFFFFFFFFFF; assign b = 64'h25FFFFFFFFFFFFFF;

    #10 $display("\n2**-606 * 2**-417:");
    #10 assign a = 64'h1A10000000000000; assign b = 64'h25E0000000000000;
    #10 assign a = 64'h1A1FFFFFFFFFFFFF; assign b = 64'h25EFFFFFFFFFFFFF;

    #10 $display("\n2**-605 * 2**-418:");
    #10 assign a = 64'h1A20000000000000; assign b = 64'h25D0000000000000;
    #10 assign a = 64'h1A2FFFFFFFFFFFFF; assign b = 64'h25DFFFFFFFFFFFFF;

    #10 $display("\n2**-604 * 2**-419:");
    #10 assign a = 64'h1A30000000000000; assign b = 64'h25C0000000000000;
    #10 assign a = 64'h1A3FFFFFFFFFFFFF; assign b = 64'h25CFFFFFFFFFFFFF;

    #10 $display("\n2**-603 * 2**-420:");
    #10 assign a = 64'h1A40000000000000; assign b = 64'h25B0000000000000;
    #10 assign a = 64'h1A4FFFFFFFFFFFFF; assign b = 64'h25BFFFFFFFFFFFFF;

    #10 $display("\n2**-602 * 2**-421:");
    #10 assign a = 64'h1A50000000000000; assign b = 64'h25A0000000000000;
    #10 assign a = 64'h1A5FFFFFFFFFFFFF; assign b = 64'h25AFFFFFFFFFFFFF;

    #10 $display("\n2**-601 * 2**-422:");
    #10 assign a = 64'h1A60000000000000; assign b = 64'h2590000000000000;
    #10 assign a = 64'h1A6FFFFFFFFFFFFF; assign b = 64'h259FFFFFFFFFFFFF;

    #10 $display("\n2**-600 * 2**-423:");
    #10 assign a = 64'h1A70000000000000; assign b = 64'h2580000000000000;
    #10 assign a = 64'h1A7FFFFFFFFFFFFF; assign b = 64'h258FFFFFFFFFFFFF;

    #10 $display("\n2**-599 * 2**-424:");
    #10 assign a = 64'h1A80000000000000; assign b = 64'h2570000000000000;
    #10 assign a = 64'h1A8FFFFFFFFFFFFF; assign b = 64'h257FFFFFFFFFFFFF;

    #10 $display("\n2**-598 * 2**-425:");
    #10 assign a = 64'h1A90000000000000; assign b = 64'h2560000000000000;
    #10 assign a = 64'h1A9FFFFFFFFFFFFF; assign b = 64'h256FFFFFFFFFFFFF;

    #10 $display("\n2**-597 * 2**-426:");
    #10 assign a = 64'h1AA0000000000000; assign b = 64'h2550000000000000;
    #10 assign a = 64'h1AAFFFFFFFFFFFFF; assign b = 64'h255FFFFFFFFFFFFF;

    #10 $display("\n2**-596 * 2**-427:");
    #10 assign a = 64'h1AB0000000000000; assign b = 64'h2540000000000000;
    #10 assign a = 64'h1ABFFFFFFFFFFFFF; assign b = 64'h254FFFFFFFFFFFFF;

    #10 $display("\n2**-595 * 2**-428:");
    #10 assign a = 64'h1AC0000000000000; assign b = 64'h2530000000000000;
    #10 assign a = 64'h1ACFFFFFFFFFFFFF; assign b = 64'h253FFFFFFFFFFFFF;

    #10 $display("\n2**-594 * 2**-429:");
    #10 assign a = 64'h1AD0000000000000; assign b = 64'h2520000000000000;
    #10 assign a = 64'h1ADFFFFFFFFFFFFF; assign b = 64'h252FFFFFFFFFFFFF;

    #10 $display("\n2**-593 * 2**-430:");
    #10 assign a = 64'h1AE0000000000000; assign b = 64'h2510000000000000;
    #10 assign a = 64'h1AEFFFFFFFFFFFFF; assign b = 64'h251FFFFFFFFFFFFF;

    #10 $display("\n2**-592 * 2**-431:");
    #10 assign a = 64'h1AF0000000000000; assign b = 64'h2500000000000000;
    #10 assign a = 64'h1AFFFFFFFFFFFFFF; assign b = 64'h250FFFFFFFFFFFFF;

    #10 $display("\n2**-591 * 2**-432:");
    #10 assign a = 64'h1B00000000000000; assign b = 64'h24F0000000000000;
    #10 assign a = 64'h1B0FFFFFFFFFFFFF; assign b = 64'h24FFFFFFFFFFFFFF;

    #10 $display("\n2**-590 * 2**-433:");
    #10 assign a = 64'h1B10000000000000; assign b = 64'h24E0000000000000;
    #10 assign a = 64'h1B1FFFFFFFFFFFFF; assign b = 64'h24EFFFFFFFFFFFFF;

    #10 $display("\n2**-589 * 2**-434:");
    #10 assign a = 64'h1B20000000000000; assign b = 64'h24D0000000000000;
    #10 assign a = 64'h1B2FFFFFFFFFFFFF; assign b = 64'h24DFFFFFFFFFFFFF;

    #10 $display("\n2**-588 * 2**-435:");
    #10 assign a = 64'h1B30000000000000; assign b = 64'h24C0000000000000;
    #10 assign a = 64'h1B3FFFFFFFFFFFFF; assign b = 64'h24CFFFFFFFFFFFFF;

    #10 $display("\n2**-587 * 2**-436:");
    #10 assign a = 64'h1B40000000000000; assign b = 64'h24B0000000000000;
    #10 assign a = 64'h1B4FFFFFFFFFFFFF; assign b = 64'h24BFFFFFFFFFFFFF;

    #10 $display("\n2**-586 * 2**-437:");
    #10 assign a = 64'h1B50000000000000; assign b = 64'h24A0000000000000;
    #10 assign a = 64'h1B5FFFFFFFFFFFFF; assign b = 64'h24AFFFFFFFFFFFFF;

    #10 $display("\n2**-585 * 2**-438:");
    #10 assign a = 64'h1B60000000000000; assign b = 64'h2490000000000000;
    #10 assign a = 64'h1B6FFFFFFFFFFFFF; assign b = 64'h249FFFFFFFFFFFFF;

    #10 $display("\n2**-584 * 2**-439:");
    #10 assign a = 64'h1B70000000000000; assign b = 64'h2480000000000000;
    #10 assign a = 64'h1B7FFFFFFFFFFFFF; assign b = 64'h248FFFFFFFFFFFFF;

    #10 $display("\n2**-583 * 2**-440:");
    #10 assign a = 64'h1B80000000000000; assign b = 64'h2470000000000000;
    #10 assign a = 64'h1B8FFFFFFFFFFFFF; assign b = 64'h247FFFFFFFFFFFFF;

    #10 $display("\n2**-582 * 2**-441:");
    #10 assign a = 64'h1B90000000000000; assign b = 64'h2460000000000000;
    #10 assign a = 64'h1B9FFFFFFFFFFFFF; assign b = 64'h246FFFFFFFFFFFFF;

    #10 $display("\n2**-581 * 2**-442:");
    #10 assign a = 64'h1BA0000000000000; assign b = 64'h2450000000000000;
    #10 assign a = 64'h1BAFFFFFFFFFFFFF; assign b = 64'h245FFFFFFFFFFFFF;

    #10 $display("\n2**-580 * 2**-443:");
    #10 assign a = 64'h1BB0000000000000; assign b = 64'h2440000000000000;
    #10 assign a = 64'h1BBFFFFFFFFFFFFF; assign b = 64'h244FFFFFFFFFFFFF;

    #10 $display("\n2**-579 * 2**-444:");
    #10 assign a = 64'h1BC0000000000000; assign b = 64'h2430000000000000;
    #10 assign a = 64'h1BCFFFFFFFFFFFFF; assign b = 64'h243FFFFFFFFFFFFF;

    #10 $display("\n2**-578 * 2**-445:");
    #10 assign a = 64'h1BD0000000000000; assign b = 64'h2420000000000000;
    #10 assign a = 64'h1BDFFFFFFFFFFFFF; assign b = 64'h242FFFFFFFFFFFFF;

    #10 $display("\n2**-577 * 2**-446:");
    #10 assign a = 64'h1BE0000000000000; assign b = 64'h2410000000000000;
    #10 assign a = 64'h1BEFFFFFFFFFFFFF; assign b = 64'h241FFFFFFFFFFFFF;

    #10 $display("\n2**-576 * 2**-447:");
    #10 assign a = 64'h1BF0000000000000; assign b = 64'h2400000000000000;
    #10 assign a = 64'h1BFFFFFFFFFFFFFF; assign b = 64'h240FFFFFFFFFFFFF;

    #10 $display("\n2**-575 * 2**-448:");
    #10 assign a = 64'h1C00000000000000; assign b = 64'h23F0000000000000;
    #10 assign a = 64'h1C0FFFFFFFFFFFFF; assign b = 64'h23FFFFFFFFFFFFFF;

    #10 $display("\n2**-574 * 2**-449:");
    #10 assign a = 64'h1C10000000000000; assign b = 64'h23E0000000000000;
    #10 assign a = 64'h1C1FFFFFFFFFFFFF; assign b = 64'h23EFFFFFFFFFFFFF;

    #10 $display("\n2**-573 * 2**-450:");
    #10 assign a = 64'h1C20000000000000; assign b = 64'h23D0000000000000;
    #10 assign a = 64'h1C2FFFFFFFFFFFFF; assign b = 64'h23DFFFFFFFFFFFFF;

    #10 $display("\n2**-572 * 2**-451:");
    #10 assign a = 64'h1C30000000000000; assign b = 64'h23C0000000000000;
    #10 assign a = 64'h1C3FFFFFFFFFFFFF; assign b = 64'h23CFFFFFFFFFFFFF;

    #10 $display("\n2**-571 * 2**-452:");
    #10 assign a = 64'h1C40000000000000; assign b = 64'h23B0000000000000;
    #10 assign a = 64'h1C4FFFFFFFFFFFFF; assign b = 64'h23BFFFFFFFFFFFFF;

    #10 $display("\n2**-570 * 2**-453:");
    #10 assign a = 64'h1C50000000000000; assign b = 64'h23A0000000000000;
    #10 assign a = 64'h1C5FFFFFFFFFFFFF; assign b = 64'h23AFFFFFFFFFFFFF;

    #10 $display("\n2**-569 * 2**-454:");
    #10 assign a = 64'h1C60000000000000; assign b = 64'h2390000000000000;
    #10 assign a = 64'h1C6FFFFFFFFFFFFF; assign b = 64'h239FFFFFFFFFFFFF;

    #10 $display("\n2**-568 * 2**-455:");
    #10 assign a = 64'h1C70000000000000; assign b = 64'h2380000000000000;
    #10 assign a = 64'h1C7FFFFFFFFFFFFF; assign b = 64'h238FFFFFFFFFFFFF;

    #10 $display("\n2**-567 * 2**-456:");
    #10 assign a = 64'h1C80000000000000; assign b = 64'h2370000000000000;
    #10 assign a = 64'h1C8FFFFFFFFFFFFF; assign b = 64'h237FFFFFFFFFFFFF;

    #10 $display("\n2**-566 * 2**-457:");
    #10 assign a = 64'h1C90000000000000; assign b = 64'h2360000000000000;
    #10 assign a = 64'h1C9FFFFFFFFFFFFF; assign b = 64'h236FFFFFFFFFFFFF;

    #10 $display("\n2**-565 * 2**-458:");
    #10 assign a = 64'h1CA0000000000000; assign b = 64'h2350000000000000;
    #10 assign a = 64'h1CAFFFFFFFFFFFFF; assign b = 64'h235FFFFFFFFFFFFF;

    #10 $display("\n2**-564 * 2**-459:");
    #10 assign a = 64'h1CB0000000000000; assign b = 64'h2340000000000000;
    #10 assign a = 64'h1CBFFFFFFFFFFFFF; assign b = 64'h234FFFFFFFFFFFFF;

    #10 $display("\n2**-563 * 2**-460:");
    #10 assign a = 64'h1CC0000000000000; assign b = 64'h2330000000000000;
    #10 assign a = 64'h1CCFFFFFFFFFFFFF; assign b = 64'h233FFFFFFFFFFFFF;

    #10 $display("\n2**-562 * 2**-461:");
    #10 assign a = 64'h1CD0000000000000; assign b = 64'h2320000000000000;
    #10 assign a = 64'h1CDFFFFFFFFFFFFF; assign b = 64'h232FFFFFFFFFFFFF;

    #10 $display("\n2**-561 * 2**-462:");
    #10 assign a = 64'h1CE0000000000000; assign b = 64'h2310000000000000;
    #10 assign a = 64'h1CEFFFFFFFFFFFFF; assign b = 64'h231FFFFFFFFFFFFF;

    #10 $display("\n2**-560 * 2**-463:");
    #10 assign a = 64'h1CF0000000000000; assign b = 64'h2300000000000000;
    #10 assign a = 64'h1CFFFFFFFFFFFFFF; assign b = 64'h230FFFFFFFFFFFFF;

    #10 $display("\n2**-559 * 2**-464:");
    #10 assign a = 64'h1D00000000000000; assign b = 64'h22F0000000000000;
    #10 assign a = 64'h1D0FFFFFFFFFFFFF; assign b = 64'h22FFFFFFFFFFFFFF;

    #10 $display("\n2**-558 * 2**-465:");
    #10 assign a = 64'h1D10000000000000; assign b = 64'h22E0000000000000;
    #10 assign a = 64'h1D1FFFFFFFFFFFFF; assign b = 64'h22EFFFFFFFFFFFFF;

    #10 $display("\n2**-557 * 2**-466:");
    #10 assign a = 64'h1D20000000000000; assign b = 64'h22D0000000000000;
    #10 assign a = 64'h1D2FFFFFFFFFFFFF; assign b = 64'h22DFFFFFFFFFFFFF;

    #10 $display("\n2**-556 * 2**-467:");
    #10 assign a = 64'h1D30000000000000; assign b = 64'h22C0000000000000;
    #10 assign a = 64'h1D3FFFFFFFFFFFFF; assign b = 64'h22CFFFFFFFFFFFFF;

    #10 $display("\n2**-555 * 2**-468:");
    #10 assign a = 64'h1D40000000000000; assign b = 64'h22B0000000000000;
    #10 assign a = 64'h1D4FFFFFFFFFFFFF; assign b = 64'h22BFFFFFFFFFFFFF;

    #10 $display("\n2**-554 * 2**-469:");
    #10 assign a = 64'h1D50000000000000; assign b = 64'h22A0000000000000;
    #10 assign a = 64'h1D5FFFFFFFFFFFFF; assign b = 64'h22AFFFFFFFFFFFFF;

    #10 $display("\n2**-553 * 2**-470:");
    #10 assign a = 64'h1D60000000000000; assign b = 64'h2290000000000000;
    #10 assign a = 64'h1D6FFFFFFFFFFFFF; assign b = 64'h229FFFFFFFFFFFFF;

    #10 $display("\n2**-552 * 2**-471:");
    #10 assign a = 64'h1D70000000000000; assign b = 64'h2280000000000000;
    #10 assign a = 64'h1D7FFFFFFFFFFFFF; assign b = 64'h228FFFFFFFFFFFFF;

    #10 $display("\n2**-551 * 2**-472:");
    #10 assign a = 64'h1D80000000000000; assign b = 64'h2270000000000000;
    #10 assign a = 64'h1D8FFFFFFFFFFFFF; assign b = 64'h227FFFFFFFFFFFFF;

    #10 $display("\n2**-550 * 2**-473:");
    #10 assign a = 64'h1D90000000000000; assign b = 64'h2260000000000000;
    #10 assign a = 64'h1D9FFFFFFFFFFFFF; assign b = 64'h226FFFFFFFFFFFFF;

    #10 $display("\n2**-549 * 2**-474:");
    #10 assign a = 64'h1DA0000000000000; assign b = 64'h2250000000000000;
    #10 assign a = 64'h1DAFFFFFFFFFFFFF; assign b = 64'h225FFFFFFFFFFFFF;

    #10 $display("\n2**-548 * 2**-475:");
    #10 assign a = 64'h1DB0000000000000; assign b = 64'h2240000000000000;
    #10 assign a = 64'h1DBFFFFFFFFFFFFF; assign b = 64'h224FFFFFFFFFFFFF;

    #10 $display("\n2**-547 * 2**-476:");
    #10 assign a = 64'h1DC0000000000000; assign b = 64'h2230000000000000;
    #10 assign a = 64'h1DCFFFFFFFFFFFFF; assign b = 64'h223FFFFFFFFFFFFF;

    #10 $display("\n2**-546 * 2**-477:");
    #10 assign a = 64'h1DD0000000000000; assign b = 64'h2220000000000000;
    #10 assign a = 64'h1DDFFFFFFFFFFFFF; assign b = 64'h222FFFFFFFFFFFFF;

    #10 $display("\n2**-545 * 2**-478:");
    #10 assign a = 64'h1DE0000000000000; assign b = 64'h2210000000000000;
    #10 assign a = 64'h1DEFFFFFFFFFFFFF; assign b = 64'h221FFFFFFFFFFFFF;

    #10 $display("\n2**-544 * 2**-479:");
    #10 assign a = 64'h1DF0000000000000; assign b = 64'h2200000000000000;
    #10 assign a = 64'h1DFFFFFFFFFFFFFF; assign b = 64'h220FFFFFFFFFFFFF;

    #10 $display("\n2**-543 * 2**-480:");
    #10 assign a = 64'h1E00000000000000; assign b = 64'h21F0000000000000;
    #10 assign a = 64'h1E0FFFFFFFFFFFFF; assign b = 64'h21FFFFFFFFFFFFFF;

    #10 $display("\n2**-542 * 2**-481:");
    #10 assign a = 64'h1E10000000000000; assign b = 64'h21E0000000000000;
    #10 assign a = 64'h1E1FFFFFFFFFFFFF; assign b = 64'h21EFFFFFFFFFFFFF;

    #10 $display("\n2**-541 * 2**-482:");
    #10 assign a = 64'h1E20000000000000; assign b = 64'h21D0000000000000;
    #10 assign a = 64'h1E2FFFFFFFFFFFFF; assign b = 64'h21DFFFFFFFFFFFFF;

    #10 $display("\n2**-540 * 2**-483:");
    #10 assign a = 64'h1E30000000000000; assign b = 64'h21C0000000000000;
    #10 assign a = 64'h1E3FFFFFFFFFFFFF; assign b = 64'h21CFFFFFFFFFFFFF;

    #10 $display("\n2**-539 * 2**-484:");
    #10 assign a = 64'h1E40000000000000; assign b = 64'h21B0000000000000;
    #10 assign a = 64'h1E4FFFFFFFFFFFFF; assign b = 64'h21BFFFFFFFFFFFFF;

    #10 $display("\n2**-538 * 2**-485:");
    #10 assign a = 64'h1E50000000000000; assign b = 64'h21A0000000000000;
    #10 assign a = 64'h1E5FFFFFFFFFFFFF; assign b = 64'h21AFFFFFFFFFFFFF;

    #10 $display("\n2**-537 * 2**-486:");
    #10 assign a = 64'h1E60000000000000; assign b = 64'h2190000000000000;
    #10 assign a = 64'h1E6FFFFFFFFFFFFF; assign b = 64'h219FFFFFFFFFFFFF;

    #10 $display("\n2**-536 * 2**-487:");
    #10 assign a = 64'h1E70000000000000; assign b = 64'h2180000000000000;
    #10 assign a = 64'h1E7FFFFFFFFFFFFF; assign b = 64'h218FFFFFFFFFFFFF;

    #10 $display("\n2**-535 * 2**-488:");
    #10 assign a = 64'h1E80000000000000; assign b = 64'h2170000000000000;
    #10 assign a = 64'h1E8FFFFFFFFFFFFF; assign b = 64'h217FFFFFFFFFFFFF;

    #10 $display("\n2**-534 * 2**-489:");
    #10 assign a = 64'h1E90000000000000; assign b = 64'h2160000000000000;
    #10 assign a = 64'h1E9FFFFFFFFFFFFF; assign b = 64'h216FFFFFFFFFFFFF;

    #10 $display("\n2**-533 * 2**-490:");
    #10 assign a = 64'h1EA0000000000000; assign b = 64'h2150000000000000;
    #10 assign a = 64'h1EAFFFFFFFFFFFFF; assign b = 64'h215FFFFFFFFFFFFF;

    #10 $display("\n2**-532 * 2**-491:");
    #10 assign a = 64'h1EB0000000000000; assign b = 64'h2140000000000000;
    #10 assign a = 64'h1EBFFFFFFFFFFFFF; assign b = 64'h214FFFFFFFFFFFFF;

    #10 $display("\n2**-531 * 2**-492:");
    #10 assign a = 64'h1EC0000000000000; assign b = 64'h2130000000000000;
    #10 assign a = 64'h1ECFFFFFFFFFFFFF; assign b = 64'h213FFFFFFFFFFFFF;

    #10 $display("\n2**-530 * 2**-493:");
    #10 assign a = 64'h1ED0000000000000; assign b = 64'h2120000000000000;
    #10 assign a = 64'h1EDFFFFFFFFFFFFF; assign b = 64'h212FFFFFFFFFFFFF;

    #10 $display("\n2**-529 * 2**-494:");
    #10 assign a = 64'h1EE0000000000000; assign b = 64'h2110000000000000;
    #10 assign a = 64'h1EEFFFFFFFFFFFFF; assign b = 64'h211FFFFFFFFFFFFF;

    #10 $display("\n2**-528 * 2**-495:");
    #10 assign a = 64'h1EF0000000000000; assign b = 64'h2100000000000000;
    #10 assign a = 64'h1EFFFFFFFFFFFFFF; assign b = 64'h210FFFFFFFFFFFFF;

    #10 $display("\n2**-527 * 2**-496:");
    #10 assign a = 64'h1F00000000000000; assign b = 64'h20F0000000000000;
    #10 assign a = 64'h1F0FFFFFFFFFFFFF; assign b = 64'h20FFFFFFFFFFFFFF;

    #10 $display("\n2**-526 * 2**-497:");
    #10 assign a = 64'h1F10000000000000; assign b = 64'h20E0000000000000;
    #10 assign a = 64'h1F1FFFFFFFFFFFFF; assign b = 64'h20EFFFFFFFFFFFFF;

    #10 $display("\n2**-525 * 2**-498:");
    #10 assign a = 64'h1F20000000000000; assign b = 64'h20D0000000000000;
    #10 assign a = 64'h1F2FFFFFFFFFFFFF; assign b = 64'h20DFFFFFFFFFFFFF;

    #10 $display("\n2**-524 * 2**-499:");
    #10 assign a = 64'h1F30000000000000; assign b = 64'h20C0000000000000;
    #10 assign a = 64'h1F3FFFFFFFFFFFFF; assign b = 64'h20CFFFFFFFFFFFFF;

    #10 $display("\n2**-523 * 2**-500:");
    #10 assign a = 64'h1F40000000000000; assign b = 64'h20B0000000000000;
    #10 assign a = 64'h1F4FFFFFFFFFFFFF; assign b = 64'h20BFFFFFFFFFFFFF;

    #10 $display("\n2**-522 * 2**-501:");
    #10 assign a = 64'h1F50000000000000; assign b = 64'h20A0000000000000;
    #10 assign a = 64'h1F5FFFFFFFFFFFFF; assign b = 64'h20AFFFFFFFFFFFFF;

    #10 $display("\n2**-521 * 2**-502:");
    #10 assign a = 64'h1F60000000000000; assign b = 64'h2090000000000000;
    #10 assign a = 64'h1F6FFFFFFFFFFFFF; assign b = 64'h209FFFFFFFFFFFFF;

    #10 $display("\n2**-520 * 2**-503:");
    #10 assign a = 64'h1F70000000000000; assign b = 64'h2080000000000000;
    #10 assign a = 64'h1F7FFFFFFFFFFFFF; assign b = 64'h208FFFFFFFFFFFFF;

    #10 $display("\n2**-519 * 2**-504:");
    #10 assign a = 64'h1F80000000000000; assign b = 64'h2070000000000000;
    #10 assign a = 64'h1F8FFFFFFFFFFFFF; assign b = 64'h207FFFFFFFFFFFFF;

    #10 $display("\n2**-518 * 2**-505:");
    #10 assign a = 64'h1F90000000000000; assign b = 64'h2060000000000000;
    #10 assign a = 64'h1F9FFFFFFFFFFFFF; assign b = 64'h206FFFFFFFFFFFFF;

    #10 $display("\n2**-517 * 2**-506:");
    #10 assign a = 64'h1FA0000000000000; assign b = 64'h2050000000000000;
    #10 assign a = 64'h1FAFFFFFFFFFFFFF; assign b = 64'h205FFFFFFFFFFFFF;

    #10 $display("\n2**-516 * 2**-507:");
    #10 assign a = 64'h1FB0000000000000; assign b = 64'h2040000000000000;
    #10 assign a = 64'h1FBFFFFFFFFFFFFF; assign b = 64'h204FFFFFFFFFFFFF;

    #10 $display("\n2**-515 * 2**-508:");
    #10 assign a = 64'h1FC0000000000000; assign b = 64'h2030000000000000;
    #10 assign a = 64'h1FCFFFFFFFFFFFFF; assign b = 64'h203FFFFFFFFFFFFF;

    #10 $display("\n2**-514 * 2**-509:");
    #10 assign a = 64'h1FD0000000000000; assign b = 64'h2020000000000000;
    #10 assign a = 64'h1FDFFFFFFFFFFFFF; assign b = 64'h202FFFFFFFFFFFFF;

    #10 $display("\n2**-513 * 2**-510:");
    #10 assign a = 64'h1FE0000000000000; assign b = 64'h2010000000000000;
    #10 assign a = 64'h1FEFFFFFFFFFFFFF; assign b = 64'h201FFFFFFFFFFFFF;

    #10 $display("\n2**-512 * 2**-511:");
    #10 assign a = 64'h1FF0000000000000; assign b = 64'h2000000000000000;
    #10 assign a = 64'h1FFFFFFFFFFFFFFF; assign b = 64'h200FFFFFFFFFFFFF;

    #10 $display("\n2**-511 * 2**-512:");
    #10 assign a = 64'h2000000000000000; assign b = 64'h1FF0000000000000;
    #10 assign a = 64'h200FFFFFFFFFFFFF; assign b = 64'h1FFFFFFFFFFFFFFF;

    #10 $display("\n2**-510 * 2**-513:");
    #10 assign a = 64'h2010000000000000; assign b = 64'h1FE0000000000000;
    #10 assign a = 64'h201FFFFFFFFFFFFF; assign b = 64'h1FEFFFFFFFFFFFFF;

    #10 $display("\n2**-509 * 2**-514:");
    #10 assign a = 64'h2020000000000000; assign b = 64'h1FD0000000000000;
    #10 assign a = 64'h202FFFFFFFFFFFFF; assign b = 64'h1FDFFFFFFFFFFFFF;

    #10 $display("\n2**-508 * 2**-515:");
    #10 assign a = 64'h2030000000000000; assign b = 64'h1FC0000000000000;
    #10 assign a = 64'h203FFFFFFFFFFFFF; assign b = 64'h1FCFFFFFFFFFFFFF;

    #10 $display("\n2**-507 * 2**-516:");
    #10 assign a = 64'h2040000000000000; assign b = 64'h1FB0000000000000;
    #10 assign a = 64'h204FFFFFFFFFFFFF; assign b = 64'h1FBFFFFFFFFFFFFF;

    #10 $display("\n2**-506 * 2**-517:");
    #10 assign a = 64'h2050000000000000; assign b = 64'h1FA0000000000000;
    #10 assign a = 64'h205FFFFFFFFFFFFF; assign b = 64'h1FAFFFFFFFFFFFFF;

    #10 $display("\n2**-505 * 2**-518:");
    #10 assign a = 64'h2060000000000000; assign b = 64'h1F90000000000000;
    #10 assign a = 64'h206FFFFFFFFFFFFF; assign b = 64'h1F9FFFFFFFFFFFFF;

    #10 $display("\n2**-504 * 2**-519:");
    #10 assign a = 64'h2070000000000000; assign b = 64'h1F80000000000000;
    #10 assign a = 64'h207FFFFFFFFFFFFF; assign b = 64'h1F8FFFFFFFFFFFFF;

    #10 $display("\n2**-503 * 2**-520:");
    #10 assign a = 64'h2080000000000000; assign b = 64'h1F70000000000000;
    #10 assign a = 64'h208FFFFFFFFFFFFF; assign b = 64'h1F7FFFFFFFFFFFFF;

    #10 $display("\n2**-502 * 2**-521:");
    #10 assign a = 64'h2090000000000000; assign b = 64'h1F60000000000000;
    #10 assign a = 64'h209FFFFFFFFFFFFF; assign b = 64'h1F6FFFFFFFFFFFFF;

    #10 $display("\n2**-501 * 2**-522:");
    #10 assign a = 64'h20A0000000000000; assign b = 64'h1F50000000000000;
    #10 assign a = 64'h20AFFFFFFFFFFFFF; assign b = 64'h1F5FFFFFFFFFFFFF;

    #10 $display("\n2**-500 * 2**-523:");
    #10 assign a = 64'h20B0000000000000; assign b = 64'h1F40000000000000;
    #10 assign a = 64'h20BFFFFFFFFFFFFF; assign b = 64'h1F4FFFFFFFFFFFFF;

    #10 $display("\n2**-499 * 2**-524:");
    #10 assign a = 64'h20C0000000000000; assign b = 64'h1F30000000000000;
    #10 assign a = 64'h20CFFFFFFFFFFFFF; assign b = 64'h1F3FFFFFFFFFFFFF;

    #10 $display("\n2**-498 * 2**-525:");
    #10 assign a = 64'h20D0000000000000; assign b = 64'h1F20000000000000;
    #10 assign a = 64'h20DFFFFFFFFFFFFF; assign b = 64'h1F2FFFFFFFFFFFFF;

    #10 $display("\n2**-497 * 2**-526:");
    #10 assign a = 64'h20E0000000000000; assign b = 64'h1F10000000000000;
    #10 assign a = 64'h20EFFFFFFFFFFFFF; assign b = 64'h1F1FFFFFFFFFFFFF;

    #10 $display("\n2**-496 * 2**-527:");
    #10 assign a = 64'h20F0000000000000; assign b = 64'h1F00000000000000;
    #10 assign a = 64'h20FFFFFFFFFFFFFF; assign b = 64'h1F0FFFFFFFFFFFFF;

    #10 $display("\n2**-495 * 2**-528:");
    #10 assign a = 64'h2100000000000000; assign b = 64'h1EF0000000000000;
    #10 assign a = 64'h210FFFFFFFFFFFFF; assign b = 64'h1EFFFFFFFFFFFFFF;

    #10 $display("\n2**-494 * 2**-529:");
    #10 assign a = 64'h2110000000000000; assign b = 64'h1EE0000000000000;
    #10 assign a = 64'h211FFFFFFFFFFFFF; assign b = 64'h1EEFFFFFFFFFFFFF;

    #10 $display("\n2**-493 * 2**-530:");
    #10 assign a = 64'h2120000000000000; assign b = 64'h1ED0000000000000;
    #10 assign a = 64'h212FFFFFFFFFFFFF; assign b = 64'h1EDFFFFFFFFFFFFF;

    #10 $display("\n2**-492 * 2**-531:");
    #10 assign a = 64'h2130000000000000; assign b = 64'h1EC0000000000000;
    #10 assign a = 64'h213FFFFFFFFFFFFF; assign b = 64'h1ECFFFFFFFFFFFFF;

    #10 $display("\n2**-491 * 2**-532:");
    #10 assign a = 64'h2140000000000000; assign b = 64'h1EB0000000000000;
    #10 assign a = 64'h214FFFFFFFFFFFFF; assign b = 64'h1EBFFFFFFFFFFFFF;

    #10 $display("\n2**-490 * 2**-533:");
    #10 assign a = 64'h2150000000000000; assign b = 64'h1EA0000000000000;
    #10 assign a = 64'h215FFFFFFFFFFFFF; assign b = 64'h1EAFFFFFFFFFFFFF;

    #10 $display("\n2**-489 * 2**-534:");
    #10 assign a = 64'h2160000000000000; assign b = 64'h1E90000000000000;
    #10 assign a = 64'h216FFFFFFFFFFFFF; assign b = 64'h1E9FFFFFFFFFFFFF;

    #10 $display("\n2**-488 * 2**-535:");
    #10 assign a = 64'h2170000000000000; assign b = 64'h1E80000000000000;
    #10 assign a = 64'h217FFFFFFFFFFFFF; assign b = 64'h1E8FFFFFFFFFFFFF;

    #10 $display("\n2**-487 * 2**-536:");
    #10 assign a = 64'h2180000000000000; assign b = 64'h1E70000000000000;
    #10 assign a = 64'h218FFFFFFFFFFFFF; assign b = 64'h1E7FFFFFFFFFFFFF;

    #10 $display("\n2**-486 * 2**-537:");
    #10 assign a = 64'h2190000000000000; assign b = 64'h1E60000000000000;
    #10 assign a = 64'h219FFFFFFFFFFFFF; assign b = 64'h1E6FFFFFFFFFFFFF;

    #10 $display("\n2**-485 * 2**-538:");
    #10 assign a = 64'h21A0000000000000; assign b = 64'h1E50000000000000;
    #10 assign a = 64'h21AFFFFFFFFFFFFF; assign b = 64'h1E5FFFFFFFFFFFFF;

    #10 $display("\n2**-484 * 2**-539:");
    #10 assign a = 64'h21B0000000000000; assign b = 64'h1E40000000000000;
    #10 assign a = 64'h21BFFFFFFFFFFFFF; assign b = 64'h1E4FFFFFFFFFFFFF;

    #10 $display("\n2**-483 * 2**-540:");
    #10 assign a = 64'h21C0000000000000; assign b = 64'h1E30000000000000;
    #10 assign a = 64'h21CFFFFFFFFFFFFF; assign b = 64'h1E3FFFFFFFFFFFFF;

    #10 $display("\n2**-482 * 2**-541:");
    #10 assign a = 64'h21D0000000000000; assign b = 64'h1E20000000000000;
    #10 assign a = 64'h21DFFFFFFFFFFFFF; assign b = 64'h1E2FFFFFFFFFFFFF;

    #10 $display("\n2**-481 * 2**-542:");
    #10 assign a = 64'h21E0000000000000; assign b = 64'h1E10000000000000;
    #10 assign a = 64'h21EFFFFFFFFFFFFF; assign b = 64'h1E1FFFFFFFFFFFFF;

    #10 $display("\n2**-480 * 2**-543:");
    #10 assign a = 64'h21F0000000000000; assign b = 64'h1E00000000000000;
    #10 assign a = 64'h21FFFFFFFFFFFFFF; assign b = 64'h1E0FFFFFFFFFFFFF;

    #10 $display("\n2**-479 * 2**-544:");
    #10 assign a = 64'h2200000000000000; assign b = 64'h1DF0000000000000;
    #10 assign a = 64'h220FFFFFFFFFFFFF; assign b = 64'h1DFFFFFFFFFFFFFF;

    #10 $display("\n2**-478 * 2**-545:");
    #10 assign a = 64'h2210000000000000; assign b = 64'h1DE0000000000000;
    #10 assign a = 64'h221FFFFFFFFFFFFF; assign b = 64'h1DEFFFFFFFFFFFFF;

    #10 $display("\n2**-477 * 2**-546:");
    #10 assign a = 64'h2220000000000000; assign b = 64'h1DD0000000000000;
    #10 assign a = 64'h222FFFFFFFFFFFFF; assign b = 64'h1DDFFFFFFFFFFFFF;

    #10 $display("\n2**-476 * 2**-547:");
    #10 assign a = 64'h2230000000000000; assign b = 64'h1DC0000000000000;
    #10 assign a = 64'h223FFFFFFFFFFFFF; assign b = 64'h1DCFFFFFFFFFFFFF;

    #10 $display("\n2**-475 * 2**-548:");
    #10 assign a = 64'h2240000000000000; assign b = 64'h1DB0000000000000;
    #10 assign a = 64'h224FFFFFFFFFFFFF; assign b = 64'h1DBFFFFFFFFFFFFF;

    #10 $display("\n2**-474 * 2**-549:");
    #10 assign a = 64'h2250000000000000; assign b = 64'h1DA0000000000000;
    #10 assign a = 64'h225FFFFFFFFFFFFF; assign b = 64'h1DAFFFFFFFFFFFFF;

    #10 $display("\n2**-473 * 2**-550:");
    #10 assign a = 64'h2260000000000000; assign b = 64'h1D90000000000000;
    #10 assign a = 64'h226FFFFFFFFFFFFF; assign b = 64'h1D9FFFFFFFFFFFFF;

    #10 $display("\n2**-472 * 2**-551:");
    #10 assign a = 64'h2270000000000000; assign b = 64'h1D80000000000000;
    #10 assign a = 64'h227FFFFFFFFFFFFF; assign b = 64'h1D8FFFFFFFFFFFFF;

    #10 $display("\n2**-471 * 2**-552:");
    #10 assign a = 64'h2280000000000000; assign b = 64'h1D70000000000000;
    #10 assign a = 64'h228FFFFFFFFFFFFF; assign b = 64'h1D7FFFFFFFFFFFFF;

    #10 $display("\n2**-470 * 2**-553:");
    #10 assign a = 64'h2290000000000000; assign b = 64'h1D60000000000000;
    #10 assign a = 64'h229FFFFFFFFFFFFF; assign b = 64'h1D6FFFFFFFFFFFFF;

    #10 $display("\n2**-469 * 2**-554:");
    #10 assign a = 64'h22A0000000000000; assign b = 64'h1D50000000000000;
    #10 assign a = 64'h22AFFFFFFFFFFFFF; assign b = 64'h1D5FFFFFFFFFFFFF;

    #10 $display("\n2**-468 * 2**-555:");
    #10 assign a = 64'h22B0000000000000; assign b = 64'h1D40000000000000;
    #10 assign a = 64'h22BFFFFFFFFFFFFF; assign b = 64'h1D4FFFFFFFFFFFFF;

    #10 $display("\n2**-467 * 2**-556:");
    #10 assign a = 64'h22C0000000000000; assign b = 64'h1D30000000000000;
    #10 assign a = 64'h22CFFFFFFFFFFFFF; assign b = 64'h1D3FFFFFFFFFFFFF;

    #10 $display("\n2**-466 * 2**-557:");
    #10 assign a = 64'h22D0000000000000; assign b = 64'h1D20000000000000;
    #10 assign a = 64'h22DFFFFFFFFFFFFF; assign b = 64'h1D2FFFFFFFFFFFFF;

    #10 $display("\n2**-465 * 2**-558:");
    #10 assign a = 64'h22E0000000000000; assign b = 64'h1D10000000000000;
    #10 assign a = 64'h22EFFFFFFFFFFFFF; assign b = 64'h1D1FFFFFFFFFFFFF;

    #10 $display("\n2**-464 * 2**-559:");
    #10 assign a = 64'h22F0000000000000; assign b = 64'h1D00000000000000;
    #10 assign a = 64'h22FFFFFFFFFFFFFF; assign b = 64'h1D0FFFFFFFFFFFFF;

    #10 $display("\n2**-463 * 2**-560:");
    #10 assign a = 64'h2300000000000000; assign b = 64'h1CF0000000000000;
    #10 assign a = 64'h230FFFFFFFFFFFFF; assign b = 64'h1CFFFFFFFFFFFFFF;

    #10 $display("\n2**-462 * 2**-561:");
    #10 assign a = 64'h2310000000000000; assign b = 64'h1CE0000000000000;
    #10 assign a = 64'h231FFFFFFFFFFFFF; assign b = 64'h1CEFFFFFFFFFFFFF;

    #10 $display("\n2**-461 * 2**-562:");
    #10 assign a = 64'h2320000000000000; assign b = 64'h1CD0000000000000;
    #10 assign a = 64'h232FFFFFFFFFFFFF; assign b = 64'h1CDFFFFFFFFFFFFF;

    #10 $display("\n2**-460 * 2**-563:");
    #10 assign a = 64'h2330000000000000; assign b = 64'h1CC0000000000000;
    #10 assign a = 64'h233FFFFFFFFFFFFF; assign b = 64'h1CCFFFFFFFFFFFFF;

    #10 $display("\n2**-459 * 2**-564:");
    #10 assign a = 64'h2340000000000000; assign b = 64'h1CB0000000000000;
    #10 assign a = 64'h234FFFFFFFFFFFFF; assign b = 64'h1CBFFFFFFFFFFFFF;

    #10 $display("\n2**-458 * 2**-565:");
    #10 assign a = 64'h2350000000000000; assign b = 64'h1CA0000000000000;
    #10 assign a = 64'h235FFFFFFFFFFFFF; assign b = 64'h1CAFFFFFFFFFFFFF;

    #10 $display("\n2**-457 * 2**-566:");
    #10 assign a = 64'h2360000000000000; assign b = 64'h1C90000000000000;
    #10 assign a = 64'h236FFFFFFFFFFFFF; assign b = 64'h1C9FFFFFFFFFFFFF;

    #10 $display("\n2**-456 * 2**-567:");
    #10 assign a = 64'h2370000000000000; assign b = 64'h1C80000000000000;
    #10 assign a = 64'h237FFFFFFFFFFFFF; assign b = 64'h1C8FFFFFFFFFFFFF;

    #10 $display("\n2**-455 * 2**-568:");
    #10 assign a = 64'h2380000000000000; assign b = 64'h1C70000000000000;
    #10 assign a = 64'h238FFFFFFFFFFFFF; assign b = 64'h1C7FFFFFFFFFFFFF;

    #10 $display("\n2**-454 * 2**-569:");
    #10 assign a = 64'h2390000000000000; assign b = 64'h1C60000000000000;
    #10 assign a = 64'h239FFFFFFFFFFFFF; assign b = 64'h1C6FFFFFFFFFFFFF;

    #10 $display("\n2**-453 * 2**-570:");
    #10 assign a = 64'h23A0000000000000; assign b = 64'h1C50000000000000;
    #10 assign a = 64'h23AFFFFFFFFFFFFF; assign b = 64'h1C5FFFFFFFFFFFFF;

    #10 $display("\n2**-452 * 2**-571:");
    #10 assign a = 64'h23B0000000000000; assign b = 64'h1C40000000000000;
    #10 assign a = 64'h23BFFFFFFFFFFFFF; assign b = 64'h1C4FFFFFFFFFFFFF;

    #10 $display("\n2**-451 * 2**-572:");
    #10 assign a = 64'h23C0000000000000; assign b = 64'h1C30000000000000;
    #10 assign a = 64'h23CFFFFFFFFFFFFF; assign b = 64'h1C3FFFFFFFFFFFFF;

    #10 $display("\n2**-450 * 2**-573:");
    #10 assign a = 64'h23D0000000000000; assign b = 64'h1C20000000000000;
    #10 assign a = 64'h23DFFFFFFFFFFFFF; assign b = 64'h1C2FFFFFFFFFFFFF;

    #10 $display("\n2**-449 * 2**-574:");
    #10 assign a = 64'h23E0000000000000; assign b = 64'h1C10000000000000;
    #10 assign a = 64'h23EFFFFFFFFFFFFF; assign b = 64'h1C1FFFFFFFFFFFFF;

    #10 $display("\n2**-448 * 2**-575:");
    #10 assign a = 64'h23F0000000000000; assign b = 64'h1C00000000000000;
    #10 assign a = 64'h23FFFFFFFFFFFFFF; assign b = 64'h1C0FFFFFFFFFFFFF;

    #10 $display("\n2**-447 * 2**-576:");
    #10 assign a = 64'h2400000000000000; assign b = 64'h1BF0000000000000;
    #10 assign a = 64'h240FFFFFFFFFFFFF; assign b = 64'h1BFFFFFFFFFFFFFF;

    #10 $display("\n2**-446 * 2**-577:");
    #10 assign a = 64'h2410000000000000; assign b = 64'h1BE0000000000000;
    #10 assign a = 64'h241FFFFFFFFFFFFF; assign b = 64'h1BEFFFFFFFFFFFFF;

    #10 $display("\n2**-445 * 2**-578:");
    #10 assign a = 64'h2420000000000000; assign b = 64'h1BD0000000000000;
    #10 assign a = 64'h242FFFFFFFFFFFFF; assign b = 64'h1BDFFFFFFFFFFFFF;

    #10 $display("\n2**-444 * 2**-579:");
    #10 assign a = 64'h2430000000000000; assign b = 64'h1BC0000000000000;
    #10 assign a = 64'h243FFFFFFFFFFFFF; assign b = 64'h1BCFFFFFFFFFFFFF;

    #10 $display("\n2**-443 * 2**-580:");
    #10 assign a = 64'h2440000000000000; assign b = 64'h1BB0000000000000;
    #10 assign a = 64'h244FFFFFFFFFFFFF; assign b = 64'h1BBFFFFFFFFFFFFF;

    #10 $display("\n2**-442 * 2**-581:");
    #10 assign a = 64'h2450000000000000; assign b = 64'h1BA0000000000000;
    #10 assign a = 64'h245FFFFFFFFFFFFF; assign b = 64'h1BAFFFFFFFFFFFFF;

    #10 $display("\n2**-441 * 2**-582:");
    #10 assign a = 64'h2460000000000000; assign b = 64'h1B90000000000000;
    #10 assign a = 64'h246FFFFFFFFFFFFF; assign b = 64'h1B9FFFFFFFFFFFFF;

    #10 $display("\n2**-440 * 2**-583:");
    #10 assign a = 64'h2470000000000000; assign b = 64'h1B80000000000000;
    #10 assign a = 64'h247FFFFFFFFFFFFF; assign b = 64'h1B8FFFFFFFFFFFFF;

    #10 $display("\n2**-439 * 2**-584:");
    #10 assign a = 64'h2480000000000000; assign b = 64'h1B70000000000000;
    #10 assign a = 64'h248FFFFFFFFFFFFF; assign b = 64'h1B7FFFFFFFFFFFFF;

    #10 $display("\n2**-438 * 2**-585:");
    #10 assign a = 64'h2490000000000000; assign b = 64'h1B60000000000000;
    #10 assign a = 64'h249FFFFFFFFFFFFF; assign b = 64'h1B6FFFFFFFFFFFFF;

    #10 $display("\n2**-437 * 2**-586:");
    #10 assign a = 64'h24A0000000000000; assign b = 64'h1B50000000000000;
    #10 assign a = 64'h24AFFFFFFFFFFFFF; assign b = 64'h1B5FFFFFFFFFFFFF;

    #10 $display("\n2**-436 * 2**-587:");
    #10 assign a = 64'h24B0000000000000; assign b = 64'h1B40000000000000;
    #10 assign a = 64'h24BFFFFFFFFFFFFF; assign b = 64'h1B4FFFFFFFFFFFFF;

    #10 $display("\n2**-435 * 2**-588:");
    #10 assign a = 64'h24C0000000000000; assign b = 64'h1B30000000000000;
    #10 assign a = 64'h24CFFFFFFFFFFFFF; assign b = 64'h1B3FFFFFFFFFFFFF;

    #10 $display("\n2**-434 * 2**-589:");
    #10 assign a = 64'h24D0000000000000; assign b = 64'h1B20000000000000;
    #10 assign a = 64'h24DFFFFFFFFFFFFF; assign b = 64'h1B2FFFFFFFFFFFFF;

    #10 $display("\n2**-433 * 2**-590:");
    #10 assign a = 64'h24E0000000000000; assign b = 64'h1B10000000000000;
    #10 assign a = 64'h24EFFFFFFFFFFFFF; assign b = 64'h1B1FFFFFFFFFFFFF;

    #10 $display("\n2**-432 * 2**-591:");
    #10 assign a = 64'h24F0000000000000; assign b = 64'h1B00000000000000;
    #10 assign a = 64'h24FFFFFFFFFFFFFF; assign b = 64'h1B0FFFFFFFFFFFFF;

    #10 $display("\n2**-431 * 2**-592:");
    #10 assign a = 64'h2500000000000000; assign b = 64'h1AF0000000000000;
    #10 assign a = 64'h250FFFFFFFFFFFFF; assign b = 64'h1AFFFFFFFFFFFFFF;

    #10 $display("\n2**-430 * 2**-593:");
    #10 assign a = 64'h2510000000000000; assign b = 64'h1AE0000000000000;
    #10 assign a = 64'h251FFFFFFFFFFFFF; assign b = 64'h1AEFFFFFFFFFFFFF;

    #10 $display("\n2**-429 * 2**-594:");
    #10 assign a = 64'h2520000000000000; assign b = 64'h1AD0000000000000;
    #10 assign a = 64'h252FFFFFFFFFFFFF; assign b = 64'h1ADFFFFFFFFFFFFF;

    #10 $display("\n2**-428 * 2**-595:");
    #10 assign a = 64'h2530000000000000; assign b = 64'h1AC0000000000000;
    #10 assign a = 64'h253FFFFFFFFFFFFF; assign b = 64'h1ACFFFFFFFFFFFFF;

    #10 $display("\n2**-427 * 2**-596:");
    #10 assign a = 64'h2540000000000000; assign b = 64'h1AB0000000000000;
    #10 assign a = 64'h254FFFFFFFFFFFFF; assign b = 64'h1ABFFFFFFFFFFFFF;

    #10 $display("\n2**-426 * 2**-597:");
    #10 assign a = 64'h2550000000000000; assign b = 64'h1AA0000000000000;
    #10 assign a = 64'h255FFFFFFFFFFFFF; assign b = 64'h1AAFFFFFFFFFFFFF;

    #10 $display("\n2**-425 * 2**-598:");
    #10 assign a = 64'h2560000000000000; assign b = 64'h1A90000000000000;
    #10 assign a = 64'h256FFFFFFFFFFFFF; assign b = 64'h1A9FFFFFFFFFFFFF;

    #10 $display("\n2**-424 * 2**-599:");
    #10 assign a = 64'h2570000000000000; assign b = 64'h1A80000000000000;
    #10 assign a = 64'h257FFFFFFFFFFFFF; assign b = 64'h1A8FFFFFFFFFFFFF;

    #10 $display("\n2**-423 * 2**-600:");
    #10 assign a = 64'h2580000000000000; assign b = 64'h1A70000000000000;
    #10 assign a = 64'h258FFFFFFFFFFFFF; assign b = 64'h1A7FFFFFFFFFFFFF;

    #10 $display("\n2**-422 * 2**-601:");
    #10 assign a = 64'h2590000000000000; assign b = 64'h1A60000000000000;
    #10 assign a = 64'h259FFFFFFFFFFFFF; assign b = 64'h1A6FFFFFFFFFFFFF;

    #10 $display("\n2**-421 * 2**-602:");
    #10 assign a = 64'h25A0000000000000; assign b = 64'h1A50000000000000;
    #10 assign a = 64'h25AFFFFFFFFFFFFF; assign b = 64'h1A5FFFFFFFFFFFFF;

    #10 $display("\n2**-420 * 2**-603:");
    #10 assign a = 64'h25B0000000000000; assign b = 64'h1A40000000000000;
    #10 assign a = 64'h25BFFFFFFFFFFFFF; assign b = 64'h1A4FFFFFFFFFFFFF;

    #10 $display("\n2**-419 * 2**-604:");
    #10 assign a = 64'h25C0000000000000; assign b = 64'h1A30000000000000;
    #10 assign a = 64'h25CFFFFFFFFFFFFF; assign b = 64'h1A3FFFFFFFFFFFFF;

    #10 $display("\n2**-418 * 2**-605:");
    #10 assign a = 64'h25D0000000000000; assign b = 64'h1A20000000000000;
    #10 assign a = 64'h25DFFFFFFFFFFFFF; assign b = 64'h1A2FFFFFFFFFFFFF;

    #10 $display("\n2**-417 * 2**-606:");
    #10 assign a = 64'h25E0000000000000; assign b = 64'h1A10000000000000;
    #10 assign a = 64'h25EFFFFFFFFFFFFF; assign b = 64'h1A1FFFFFFFFFFFFF;

    #10 $display("\n2**-416 * 2**-607:");
    #10 assign a = 64'h25F0000000000000; assign b = 64'h1A00000000000000;
    #10 assign a = 64'h25FFFFFFFFFFFFFF; assign b = 64'h1A0FFFFFFFFFFFFF;

    #10 $display("\n2**-415 * 2**-608:");
    #10 assign a = 64'h2600000000000000; assign b = 64'h19F0000000000000;
    #10 assign a = 64'h260FFFFFFFFFFFFF; assign b = 64'h19FFFFFFFFFFFFFF;

    #10 $display("\n2**-414 * 2**-609:");
    #10 assign a = 64'h2610000000000000; assign b = 64'h19E0000000000000;
    #10 assign a = 64'h261FFFFFFFFFFFFF; assign b = 64'h19EFFFFFFFFFFFFF;

    #10 $display("\n2**-413 * 2**-610:");
    #10 assign a = 64'h2620000000000000; assign b = 64'h19D0000000000000;
    #10 assign a = 64'h262FFFFFFFFFFFFF; assign b = 64'h19DFFFFFFFFFFFFF;

    #10 $display("\n2**-412 * 2**-611:");
    #10 assign a = 64'h2630000000000000; assign b = 64'h19C0000000000000;
    #10 assign a = 64'h263FFFFFFFFFFFFF; assign b = 64'h19CFFFFFFFFFFFFF;

    #10 $display("\n2**-411 * 2**-612:");
    #10 assign a = 64'h2640000000000000; assign b = 64'h19B0000000000000;
    #10 assign a = 64'h264FFFFFFFFFFFFF; assign b = 64'h19BFFFFFFFFFFFFF;

    #10 $display("\n2**-410 * 2**-613:");
    #10 assign a = 64'h2650000000000000; assign b = 64'h19A0000000000000;
    #10 assign a = 64'h265FFFFFFFFFFFFF; assign b = 64'h19AFFFFFFFFFFFFF;

    #10 $display("\n2**-409 * 2**-614:");
    #10 assign a = 64'h2660000000000000; assign b = 64'h1990000000000000;
    #10 assign a = 64'h266FFFFFFFFFFFFF; assign b = 64'h199FFFFFFFFFFFFF;

    #10 $display("\n2**-408 * 2**-615:");
    #10 assign a = 64'h2670000000000000; assign b = 64'h1980000000000000;
    #10 assign a = 64'h267FFFFFFFFFFFFF; assign b = 64'h198FFFFFFFFFFFFF;

    #10 $display("\n2**-407 * 2**-616:");
    #10 assign a = 64'h2680000000000000; assign b = 64'h1970000000000000;
    #10 assign a = 64'h268FFFFFFFFFFFFF; assign b = 64'h197FFFFFFFFFFFFF;

    #10 $display("\n2**-406 * 2**-617:");
    #10 assign a = 64'h2690000000000000; assign b = 64'h1960000000000000;
    #10 assign a = 64'h269FFFFFFFFFFFFF; assign b = 64'h196FFFFFFFFFFFFF;

    #10 $display("\n2**-405 * 2**-618:");
    #10 assign a = 64'h26A0000000000000; assign b = 64'h1950000000000000;
    #10 assign a = 64'h26AFFFFFFFFFFFFF; assign b = 64'h195FFFFFFFFFFFFF;

    #10 $display("\n2**-404 * 2**-619:");
    #10 assign a = 64'h26B0000000000000; assign b = 64'h1940000000000000;
    #10 assign a = 64'h26BFFFFFFFFFFFFF; assign b = 64'h194FFFFFFFFFFFFF;

    #10 $display("\n2**-403 * 2**-620:");
    #10 assign a = 64'h26C0000000000000; assign b = 64'h1930000000000000;
    #10 assign a = 64'h26CFFFFFFFFFFFFF; assign b = 64'h193FFFFFFFFFFFFF;

    #10 $display("\n2**-402 * 2**-621:");
    #10 assign a = 64'h26D0000000000000; assign b = 64'h1920000000000000;
    #10 assign a = 64'h26DFFFFFFFFFFFFF; assign b = 64'h192FFFFFFFFFFFFF;

    #10 $display("\n2**-401 * 2**-622:");
    #10 assign a = 64'h26E0000000000000; assign b = 64'h1910000000000000;
    #10 assign a = 64'h26EFFFFFFFFFFFFF; assign b = 64'h191FFFFFFFFFFFFF;

    #10 $display("\n2**-400 * 2**-623:");
    #10 assign a = 64'h26F0000000000000; assign b = 64'h1900000000000000;
    #10 assign a = 64'h26FFFFFFFFFFFFFF; assign b = 64'h190FFFFFFFFFFFFF;

    #10 $display("\n2**-399 * 2**-624:");
    #10 assign a = 64'h2700000000000000; assign b = 64'h18F0000000000000;
    #10 assign a = 64'h270FFFFFFFFFFFFF; assign b = 64'h18FFFFFFFFFFFFFF;

    #10 $display("\n2**-398 * 2**-625:");
    #10 assign a = 64'h2710000000000000; assign b = 64'h18E0000000000000;
    #10 assign a = 64'h271FFFFFFFFFFFFF; assign b = 64'h18EFFFFFFFFFFFFF;

    #10 $display("\n2**-397 * 2**-626:");
    #10 assign a = 64'h2720000000000000; assign b = 64'h18D0000000000000;
    #10 assign a = 64'h272FFFFFFFFFFFFF; assign b = 64'h18DFFFFFFFFFFFFF;

    #10 $display("\n2**-396 * 2**-627:");
    #10 assign a = 64'h2730000000000000; assign b = 64'h18C0000000000000;
    #10 assign a = 64'h273FFFFFFFFFFFFF; assign b = 64'h18CFFFFFFFFFFFFF;

    #10 $display("\n2**-395 * 2**-628:");
    #10 assign a = 64'h2740000000000000; assign b = 64'h18B0000000000000;
    #10 assign a = 64'h274FFFFFFFFFFFFF; assign b = 64'h18BFFFFFFFFFFFFF;

    #10 $display("\n2**-394 * 2**-629:");
    #10 assign a = 64'h2750000000000000; assign b = 64'h18A0000000000000;
    #10 assign a = 64'h275FFFFFFFFFFFFF; assign b = 64'h18AFFFFFFFFFFFFF;

    #10 $display("\n2**-393 * 2**-630:");
    #10 assign a = 64'h2760000000000000; assign b = 64'h1890000000000000;
    #10 assign a = 64'h276FFFFFFFFFFFFF; assign b = 64'h189FFFFFFFFFFFFF;

    #10 $display("\n2**-392 * 2**-631:");
    #10 assign a = 64'h2770000000000000; assign b = 64'h1880000000000000;
    #10 assign a = 64'h277FFFFFFFFFFFFF; assign b = 64'h188FFFFFFFFFFFFF;

    #10 $display("\n2**-391 * 2**-632:");
    #10 assign a = 64'h2780000000000000; assign b = 64'h1870000000000000;
    #10 assign a = 64'h278FFFFFFFFFFFFF; assign b = 64'h187FFFFFFFFFFFFF;

    #10 $display("\n2**-390 * 2**-633:");
    #10 assign a = 64'h2790000000000000; assign b = 64'h1860000000000000;
    #10 assign a = 64'h279FFFFFFFFFFFFF; assign b = 64'h186FFFFFFFFFFFFF;

    #10 $display("\n2**-389 * 2**-634:");
    #10 assign a = 64'h27A0000000000000; assign b = 64'h1850000000000000;
    #10 assign a = 64'h27AFFFFFFFFFFFFF; assign b = 64'h185FFFFFFFFFFFFF;

    #10 $display("\n2**-388 * 2**-635:");
    #10 assign a = 64'h27B0000000000000; assign b = 64'h1840000000000000;
    #10 assign a = 64'h27BFFFFFFFFFFFFF; assign b = 64'h184FFFFFFFFFFFFF;

    #10 $display("\n2**-387 * 2**-636:");
    #10 assign a = 64'h27C0000000000000; assign b = 64'h1830000000000000;
    #10 assign a = 64'h27CFFFFFFFFFFFFF; assign b = 64'h183FFFFFFFFFFFFF;

    #10 $display("\n2**-386 * 2**-637:");
    #10 assign a = 64'h27D0000000000000; assign b = 64'h1820000000000000;
    #10 assign a = 64'h27DFFFFFFFFFFFFF; assign b = 64'h182FFFFFFFFFFFFF;

    #10 $display("\n2**-385 * 2**-638:");
    #10 assign a = 64'h27E0000000000000; assign b = 64'h1810000000000000;
    #10 assign a = 64'h27EFFFFFFFFFFFFF; assign b = 64'h181FFFFFFFFFFFFF;

    #10 $display("\n2**-384 * 2**-639:");
    #10 assign a = 64'h27F0000000000000; assign b = 64'h1800000000000000;
    #10 assign a = 64'h27FFFFFFFFFFFFFF; assign b = 64'h180FFFFFFFFFFFFF;

    #10 $display("\n2**-383 * 2**-640:");
    #10 assign a = 64'h2800000000000000; assign b = 64'h17F0000000000000;
    #10 assign a = 64'h280FFFFFFFFFFFFF; assign b = 64'h17FFFFFFFFFFFFFF;

    #10 $display("\n2**-382 * 2**-641:");
    #10 assign a = 64'h2810000000000000; assign b = 64'h17E0000000000000;
    #10 assign a = 64'h281FFFFFFFFFFFFF; assign b = 64'h17EFFFFFFFFFFFFF;

    #10 $display("\n2**-381 * 2**-642:");
    #10 assign a = 64'h2820000000000000; assign b = 64'h17D0000000000000;
    #10 assign a = 64'h282FFFFFFFFFFFFF; assign b = 64'h17DFFFFFFFFFFFFF;

    #10 $display("\n2**-380 * 2**-643:");
    #10 assign a = 64'h2830000000000000; assign b = 64'h17C0000000000000;
    #10 assign a = 64'h283FFFFFFFFFFFFF; assign b = 64'h17CFFFFFFFFFFFFF;

    #10 $display("\n2**-379 * 2**-644:");
    #10 assign a = 64'h2840000000000000; assign b = 64'h17B0000000000000;
    #10 assign a = 64'h284FFFFFFFFFFFFF; assign b = 64'h17BFFFFFFFFFFFFF;

    #10 $display("\n2**-378 * 2**-645:");
    #10 assign a = 64'h2850000000000000; assign b = 64'h17A0000000000000;
    #10 assign a = 64'h285FFFFFFFFFFFFF; assign b = 64'h17AFFFFFFFFFFFFF;

    #10 $display("\n2**-377 * 2**-646:");
    #10 assign a = 64'h2860000000000000; assign b = 64'h1790000000000000;
    #10 assign a = 64'h286FFFFFFFFFFFFF; assign b = 64'h179FFFFFFFFFFFFF;

    #10 $display("\n2**-376 * 2**-647:");
    #10 assign a = 64'h2870000000000000; assign b = 64'h1780000000000000;
    #10 assign a = 64'h287FFFFFFFFFFFFF; assign b = 64'h178FFFFFFFFFFFFF;

    #10 $display("\n2**-375 * 2**-648:");
    #10 assign a = 64'h2880000000000000; assign b = 64'h1770000000000000;
    #10 assign a = 64'h288FFFFFFFFFFFFF; assign b = 64'h177FFFFFFFFFFFFF;

    #10 $display("\n2**-374 * 2**-649:");
    #10 assign a = 64'h2890000000000000; assign b = 64'h1760000000000000;
    #10 assign a = 64'h289FFFFFFFFFFFFF; assign b = 64'h176FFFFFFFFFFFFF;

    #10 $display("\n2**-373 * 2**-650:");
    #10 assign a = 64'h28A0000000000000; assign b = 64'h1750000000000000;
    #10 assign a = 64'h28AFFFFFFFFFFFFF; assign b = 64'h175FFFFFFFFFFFFF;

    #10 $display("\n2**-372 * 2**-651:");
    #10 assign a = 64'h28B0000000000000; assign b = 64'h1740000000000000;
    #10 assign a = 64'h28BFFFFFFFFFFFFF; assign b = 64'h174FFFFFFFFFFFFF;

    #10 $display("\n2**-371 * 2**-652:");
    #10 assign a = 64'h28C0000000000000; assign b = 64'h1730000000000000;
    #10 assign a = 64'h28CFFFFFFFFFFFFF; assign b = 64'h173FFFFFFFFFFFFF;

    #10 $display("\n2**-370 * 2**-653:");
    #10 assign a = 64'h28D0000000000000; assign b = 64'h1720000000000000;
    #10 assign a = 64'h28DFFFFFFFFFFFFF; assign b = 64'h172FFFFFFFFFFFFF;

    #10 $display("\n2**-369 * 2**-654:");
    #10 assign a = 64'h28E0000000000000; assign b = 64'h1710000000000000;
    #10 assign a = 64'h28EFFFFFFFFFFFFF; assign b = 64'h171FFFFFFFFFFFFF;

    #10 $display("\n2**-368 * 2**-655:");
    #10 assign a = 64'h28F0000000000000; assign b = 64'h1700000000000000;
    #10 assign a = 64'h28FFFFFFFFFFFFFF; assign b = 64'h170FFFFFFFFFFFFF;

    #10 $display("\n2**-367 * 2**-656:");
    #10 assign a = 64'h2900000000000000; assign b = 64'h16F0000000000000;
    #10 assign a = 64'h290FFFFFFFFFFFFF; assign b = 64'h16FFFFFFFFFFFFFF;

    #10 $display("\n2**-366 * 2**-657:");
    #10 assign a = 64'h2910000000000000; assign b = 64'h16E0000000000000;
    #10 assign a = 64'h291FFFFFFFFFFFFF; assign b = 64'h16EFFFFFFFFFFFFF;

    #10 $display("\n2**-365 * 2**-658:");
    #10 assign a = 64'h2920000000000000; assign b = 64'h16D0000000000000;
    #10 assign a = 64'h292FFFFFFFFFFFFF; assign b = 64'h16DFFFFFFFFFFFFF;

    #10 $display("\n2**-364 * 2**-659:");
    #10 assign a = 64'h2930000000000000; assign b = 64'h16C0000000000000;
    #10 assign a = 64'h293FFFFFFFFFFFFF; assign b = 64'h16CFFFFFFFFFFFFF;

    #10 $display("\n2**-363 * 2**-660:");
    #10 assign a = 64'h2940000000000000; assign b = 64'h16B0000000000000;
    #10 assign a = 64'h294FFFFFFFFFFFFF; assign b = 64'h16BFFFFFFFFFFFFF;

    #10 $display("\n2**-362 * 2**-661:");
    #10 assign a = 64'h2950000000000000; assign b = 64'h16A0000000000000;
    #10 assign a = 64'h295FFFFFFFFFFFFF; assign b = 64'h16AFFFFFFFFFFFFF;

    #10 $display("\n2**-361 * 2**-662:");
    #10 assign a = 64'h2960000000000000; assign b = 64'h1690000000000000;
    #10 assign a = 64'h296FFFFFFFFFFFFF; assign b = 64'h169FFFFFFFFFFFFF;

    #10 $display("\n2**-360 * 2**-663:");
    #10 assign a = 64'h2970000000000000; assign b = 64'h1680000000000000;
    #10 assign a = 64'h297FFFFFFFFFFFFF; assign b = 64'h168FFFFFFFFFFFFF;

    #10 $display("\n2**-359 * 2**-664:");
    #10 assign a = 64'h2980000000000000; assign b = 64'h1670000000000000;
    #10 assign a = 64'h298FFFFFFFFFFFFF; assign b = 64'h167FFFFFFFFFFFFF;

    #10 $display("\n2**-358 * 2**-665:");
    #10 assign a = 64'h2990000000000000; assign b = 64'h1660000000000000;
    #10 assign a = 64'h299FFFFFFFFFFFFF; assign b = 64'h166FFFFFFFFFFFFF;

    #10 $display("\n2**-357 * 2**-666:");
    #10 assign a = 64'h29A0000000000000; assign b = 64'h1650000000000000;
    #10 assign a = 64'h29AFFFFFFFFFFFFF; assign b = 64'h165FFFFFFFFFFFFF;

    #10 $display("\n2**-356 * 2**-667:");
    #10 assign a = 64'h29B0000000000000; assign b = 64'h1640000000000000;
    #10 assign a = 64'h29BFFFFFFFFFFFFF; assign b = 64'h164FFFFFFFFFFFFF;

    #10 $display("\n2**-355 * 2**-668:");
    #10 assign a = 64'h29C0000000000000; assign b = 64'h1630000000000000;
    #10 assign a = 64'h29CFFFFFFFFFFFFF; assign b = 64'h163FFFFFFFFFFFFF;

    #10 $display("\n2**-354 * 2**-669:");
    #10 assign a = 64'h29D0000000000000; assign b = 64'h1620000000000000;
    #10 assign a = 64'h29DFFFFFFFFFFFFF; assign b = 64'h162FFFFFFFFFFFFF;

    #10 $display("\n2**-353 * 2**-670:");
    #10 assign a = 64'h29E0000000000000; assign b = 64'h1610000000000000;
    #10 assign a = 64'h29EFFFFFFFFFFFFF; assign b = 64'h161FFFFFFFFFFFFF;

    #10 $display("\n2**-352 * 2**-671:");
    #10 assign a = 64'h29F0000000000000; assign b = 64'h1600000000000000;
    #10 assign a = 64'h29FFFFFFFFFFFFFF; assign b = 64'h160FFFFFFFFFFFFF;

    #10 $display("\n2**-351 * 2**-672:");
    #10 assign a = 64'h2A00000000000000; assign b = 64'h15F0000000000000;
    #10 assign a = 64'h2A0FFFFFFFFFFFFF; assign b = 64'h15FFFFFFFFFFFFFF;

    #10 $display("\n2**-350 * 2**-673:");
    #10 assign a = 64'h2A10000000000000; assign b = 64'h15E0000000000000;
    #10 assign a = 64'h2A1FFFFFFFFFFFFF; assign b = 64'h15EFFFFFFFFFFFFF;

    #10 $display("\n2**-349 * 2**-674:");
    #10 assign a = 64'h2A20000000000000; assign b = 64'h15D0000000000000;
    #10 assign a = 64'h2A2FFFFFFFFFFFFF; assign b = 64'h15DFFFFFFFFFFFFF;

    #10 $display("\n2**-348 * 2**-675:");
    #10 assign a = 64'h2A30000000000000; assign b = 64'h15C0000000000000;
    #10 assign a = 64'h2A3FFFFFFFFFFFFF; assign b = 64'h15CFFFFFFFFFFFFF;

    #10 $display("\n2**-347 * 2**-676:");
    #10 assign a = 64'h2A40000000000000; assign b = 64'h15B0000000000000;
    #10 assign a = 64'h2A4FFFFFFFFFFFFF; assign b = 64'h15BFFFFFFFFFFFFF;

    #10 $display("\n2**-346 * 2**-677:");
    #10 assign a = 64'h2A50000000000000; assign b = 64'h15A0000000000000;
    #10 assign a = 64'h2A5FFFFFFFFFFFFF; assign b = 64'h15AFFFFFFFFFFFFF;

    #10 $display("\n2**-345 * 2**-678:");
    #10 assign a = 64'h2A60000000000000; assign b = 64'h1590000000000000;
    #10 assign a = 64'h2A6FFFFFFFFFFFFF; assign b = 64'h159FFFFFFFFFFFFF;

    #10 $display("\n2**-344 * 2**-679:");
    #10 assign a = 64'h2A70000000000000; assign b = 64'h1580000000000000;
    #10 assign a = 64'h2A7FFFFFFFFFFFFF; assign b = 64'h158FFFFFFFFFFFFF;

    #10 $display("\n2**-343 * 2**-680:");
    #10 assign a = 64'h2A80000000000000; assign b = 64'h1570000000000000;
    #10 assign a = 64'h2A8FFFFFFFFFFFFF; assign b = 64'h157FFFFFFFFFFFFF;

    #10 $display("\n2**-342 * 2**-681:");
    #10 assign a = 64'h2A90000000000000; assign b = 64'h1560000000000000;
    #10 assign a = 64'h2A9FFFFFFFFFFFFF; assign b = 64'h156FFFFFFFFFFFFF;

    #10 $display("\n2**-341 * 2**-682:");
    #10 assign a = 64'h2AA0000000000000; assign b = 64'h1550000000000000;
    #10 assign a = 64'h2AAFFFFFFFFFFFFF; assign b = 64'h155FFFFFFFFFFFFF;

    #10 $display("\n2**-340 * 2**-683:");
    #10 assign a = 64'h2AB0000000000000; assign b = 64'h1540000000000000;
    #10 assign a = 64'h2ABFFFFFFFFFFFFF; assign b = 64'h154FFFFFFFFFFFFF;

    #10 $display("\n2**-339 * 2**-684:");
    #10 assign a = 64'h2AC0000000000000; assign b = 64'h1530000000000000;
    #10 assign a = 64'h2ACFFFFFFFFFFFFF; assign b = 64'h153FFFFFFFFFFFFF;

    #10 $display("\n2**-338 * 2**-685:");
    #10 assign a = 64'h2AD0000000000000; assign b = 64'h1520000000000000;
    #10 assign a = 64'h2ADFFFFFFFFFFFFF; assign b = 64'h152FFFFFFFFFFFFF;

    #10 $display("\n2**-337 * 2**-686:");
    #10 assign a = 64'h2AE0000000000000; assign b = 64'h1510000000000000;
    #10 assign a = 64'h2AEFFFFFFFFFFFFF; assign b = 64'h151FFFFFFFFFFFFF;

    #10 $display("\n2**-336 * 2**-687:");
    #10 assign a = 64'h2AF0000000000000; assign b = 64'h1500000000000000;
    #10 assign a = 64'h2AFFFFFFFFFFFFFF; assign b = 64'h150FFFFFFFFFFFFF;

    #10 $display("\n2**-335 * 2**-688:");
    #10 assign a = 64'h2B00000000000000; assign b = 64'h14F0000000000000;
    #10 assign a = 64'h2B0FFFFFFFFFFFFF; assign b = 64'h14FFFFFFFFFFFFFF;

    #10 $display("\n2**-334 * 2**-689:");
    #10 assign a = 64'h2B10000000000000; assign b = 64'h14E0000000000000;
    #10 assign a = 64'h2B1FFFFFFFFFFFFF; assign b = 64'h14EFFFFFFFFFFFFF;

    #10 $display("\n2**-333 * 2**-690:");
    #10 assign a = 64'h2B20000000000000; assign b = 64'h14D0000000000000;
    #10 assign a = 64'h2B2FFFFFFFFFFFFF; assign b = 64'h14DFFFFFFFFFFFFF;

    #10 $display("\n2**-332 * 2**-691:");
    #10 assign a = 64'h2B30000000000000; assign b = 64'h14C0000000000000;
    #10 assign a = 64'h2B3FFFFFFFFFFFFF; assign b = 64'h14CFFFFFFFFFFFFF;

    #10 $display("\n2**-331 * 2**-692:");
    #10 assign a = 64'h2B40000000000000; assign b = 64'h14B0000000000000;
    #10 assign a = 64'h2B4FFFFFFFFFFFFF; assign b = 64'h14BFFFFFFFFFFFFF;

    #10 $display("\n2**-330 * 2**-693:");
    #10 assign a = 64'h2B50000000000000; assign b = 64'h14A0000000000000;
    #10 assign a = 64'h2B5FFFFFFFFFFFFF; assign b = 64'h14AFFFFFFFFFFFFF;

    #10 $display("\n2**-329 * 2**-694:");
    #10 assign a = 64'h2B60000000000000; assign b = 64'h1490000000000000;
    #10 assign a = 64'h2B6FFFFFFFFFFFFF; assign b = 64'h149FFFFFFFFFFFFF;

    #10 $display("\n2**-328 * 2**-695:");
    #10 assign a = 64'h2B70000000000000; assign b = 64'h1480000000000000;
    #10 assign a = 64'h2B7FFFFFFFFFFFFF; assign b = 64'h148FFFFFFFFFFFFF;

    #10 $display("\n2**-327 * 2**-696:");
    #10 assign a = 64'h2B80000000000000; assign b = 64'h1470000000000000;
    #10 assign a = 64'h2B8FFFFFFFFFFFFF; assign b = 64'h147FFFFFFFFFFFFF;

    #10 $display("\n2**-326 * 2**-697:");
    #10 assign a = 64'h2B90000000000000; assign b = 64'h1460000000000000;
    #10 assign a = 64'h2B9FFFFFFFFFFFFF; assign b = 64'h146FFFFFFFFFFFFF;

    #10 $display("\n2**-325 * 2**-698:");
    #10 assign a = 64'h2BA0000000000000; assign b = 64'h1450000000000000;
    #10 assign a = 64'h2BAFFFFFFFFFFFFF; assign b = 64'h145FFFFFFFFFFFFF;

    #10 $display("\n2**-324 * 2**-699:");
    #10 assign a = 64'h2BB0000000000000; assign b = 64'h1440000000000000;
    #10 assign a = 64'h2BBFFFFFFFFFFFFF; assign b = 64'h144FFFFFFFFFFFFF;

    #10 $display("\n2**-323 * 2**-700:");
    #10 assign a = 64'h2BC0000000000000; assign b = 64'h1430000000000000;
    #10 assign a = 64'h2BCFFFFFFFFFFFFF; assign b = 64'h143FFFFFFFFFFFFF;

    #10 $display("\n2**-322 * 2**-701:");
    #10 assign a = 64'h2BD0000000000000; assign b = 64'h1420000000000000;
    #10 assign a = 64'h2BDFFFFFFFFFFFFF; assign b = 64'h142FFFFFFFFFFFFF;

    #10 $display("\n2**-321 * 2**-702:");
    #10 assign a = 64'h2BE0000000000000; assign b = 64'h1410000000000000;
    #10 assign a = 64'h2BEFFFFFFFFFFFFF; assign b = 64'h141FFFFFFFFFFFFF;

    #10 $display("\n2**-320 * 2**-703:");
    #10 assign a = 64'h2BF0000000000000; assign b = 64'h1400000000000000;
    #10 assign a = 64'h2BFFFFFFFFFFFFFF; assign b = 64'h140FFFFFFFFFFFFF;

    #10 $display("\n2**-319 * 2**-704:");
    #10 assign a = 64'h2C00000000000000; assign b = 64'h13F0000000000000;
    #10 assign a = 64'h2C0FFFFFFFFFFFFF; assign b = 64'h13FFFFFFFFFFFFFF;

    #10 $display("\n2**-318 * 2**-705:");
    #10 assign a = 64'h2C10000000000000; assign b = 64'h13E0000000000000;
    #10 assign a = 64'h2C1FFFFFFFFFFFFF; assign b = 64'h13EFFFFFFFFFFFFF;

    #10 $display("\n2**-317 * 2**-706:");
    #10 assign a = 64'h2C20000000000000; assign b = 64'h13D0000000000000;
    #10 assign a = 64'h2C2FFFFFFFFFFFFF; assign b = 64'h13DFFFFFFFFFFFFF;

    #10 $display("\n2**-316 * 2**-707:");
    #10 assign a = 64'h2C30000000000000; assign b = 64'h13C0000000000000;
    #10 assign a = 64'h2C3FFFFFFFFFFFFF; assign b = 64'h13CFFFFFFFFFFFFF;

    #10 $display("\n2**-315 * 2**-708:");
    #10 assign a = 64'h2C40000000000000; assign b = 64'h13B0000000000000;
    #10 assign a = 64'h2C4FFFFFFFFFFFFF; assign b = 64'h13BFFFFFFFFFFFFF;

    #10 $display("\n2**-314 * 2**-709:");
    #10 assign a = 64'h2C50000000000000; assign b = 64'h13A0000000000000;
    #10 assign a = 64'h2C5FFFFFFFFFFFFF; assign b = 64'h13AFFFFFFFFFFFFF;

    #10 $display("\n2**-313 * 2**-710:");
    #10 assign a = 64'h2C60000000000000; assign b = 64'h1390000000000000;
    #10 assign a = 64'h2C6FFFFFFFFFFFFF; assign b = 64'h139FFFFFFFFFFFFF;

    #10 $display("\n2**-312 * 2**-711:");
    #10 assign a = 64'h2C70000000000000; assign b = 64'h1380000000000000;
    #10 assign a = 64'h2C7FFFFFFFFFFFFF; assign b = 64'h138FFFFFFFFFFFFF;

    #10 $display("\n2**-311 * 2**-712:");
    #10 assign a = 64'h2C80000000000000; assign b = 64'h1370000000000000;
    #10 assign a = 64'h2C8FFFFFFFFFFFFF; assign b = 64'h137FFFFFFFFFFFFF;

    #10 $display("\n2**-310 * 2**-713:");
    #10 assign a = 64'h2C90000000000000; assign b = 64'h1360000000000000;
    #10 assign a = 64'h2C9FFFFFFFFFFFFF; assign b = 64'h136FFFFFFFFFFFFF;

    #10 $display("\n2**-309 * 2**-714:");
    #10 assign a = 64'h2CA0000000000000; assign b = 64'h1350000000000000;
    #10 assign a = 64'h2CAFFFFFFFFFFFFF; assign b = 64'h135FFFFFFFFFFFFF;

    #10 $display("\n2**-308 * 2**-715:");
    #10 assign a = 64'h2CB0000000000000; assign b = 64'h1340000000000000;
    #10 assign a = 64'h2CBFFFFFFFFFFFFF; assign b = 64'h134FFFFFFFFFFFFF;

    #10 $display("\n2**-307 * 2**-716:");
    #10 assign a = 64'h2CC0000000000000; assign b = 64'h1330000000000000;
    #10 assign a = 64'h2CCFFFFFFFFFFFFF; assign b = 64'h133FFFFFFFFFFFFF;

    #10 $display("\n2**-306 * 2**-717:");
    #10 assign a = 64'h2CD0000000000000; assign b = 64'h1320000000000000;
    #10 assign a = 64'h2CDFFFFFFFFFFFFF; assign b = 64'h132FFFFFFFFFFFFF;

    #10 $display("\n2**-305 * 2**-718:");
    #10 assign a = 64'h2CE0000000000000; assign b = 64'h1310000000000000;
    #10 assign a = 64'h2CEFFFFFFFFFFFFF; assign b = 64'h131FFFFFFFFFFFFF;

    #10 $display("\n2**-304 * 2**-719:");
    #10 assign a = 64'h2CF0000000000000; assign b = 64'h1300000000000000;
    #10 assign a = 64'h2CFFFFFFFFFFFFFF; assign b = 64'h130FFFFFFFFFFFFF;

    #10 $display("\n2**-303 * 2**-720:");
    #10 assign a = 64'h2D00000000000000; assign b = 64'h12F0000000000000;
    #10 assign a = 64'h2D0FFFFFFFFFFFFF; assign b = 64'h12FFFFFFFFFFFFFF;

    #10 $display("\n2**-302 * 2**-721:");
    #10 assign a = 64'h2D10000000000000; assign b = 64'h12E0000000000000;
    #10 assign a = 64'h2D1FFFFFFFFFFFFF; assign b = 64'h12EFFFFFFFFFFFFF;

    #10 $display("\n2**-301 * 2**-722:");
    #10 assign a = 64'h2D20000000000000; assign b = 64'h12D0000000000000;
    #10 assign a = 64'h2D2FFFFFFFFFFFFF; assign b = 64'h12DFFFFFFFFFFFFF;

    #10 $display("\n2**-300 * 2**-723:");
    #10 assign a = 64'h2D30000000000000; assign b = 64'h12C0000000000000;
    #10 assign a = 64'h2D3FFFFFFFFFFFFF; assign b = 64'h12CFFFFFFFFFFFFF;

    #10 $display("\n2**-299 * 2**-724:");
    #10 assign a = 64'h2D40000000000000; assign b = 64'h12B0000000000000;
    #10 assign a = 64'h2D4FFFFFFFFFFFFF; assign b = 64'h12BFFFFFFFFFFFFF;

    #10 $display("\n2**-298 * 2**-725:");
    #10 assign a = 64'h2D50000000000000; assign b = 64'h12A0000000000000;
    #10 assign a = 64'h2D5FFFFFFFFFFFFF; assign b = 64'h12AFFFFFFFFFFFFF;

    #10 $display("\n2**-297 * 2**-726:");
    #10 assign a = 64'h2D60000000000000; assign b = 64'h1290000000000000;
    #10 assign a = 64'h2D6FFFFFFFFFFFFF; assign b = 64'h129FFFFFFFFFFFFF;

    #10 $display("\n2**-296 * 2**-727:");
    #10 assign a = 64'h2D70000000000000; assign b = 64'h1280000000000000;
    #10 assign a = 64'h2D7FFFFFFFFFFFFF; assign b = 64'h128FFFFFFFFFFFFF;

    #10 $display("\n2**-295 * 2**-728:");
    #10 assign a = 64'h2D80000000000000; assign b = 64'h1270000000000000;
    #10 assign a = 64'h2D8FFFFFFFFFFFFF; assign b = 64'h127FFFFFFFFFFFFF;

    #10 $display("\n2**-294 * 2**-729:");
    #10 assign a = 64'h2D90000000000000; assign b = 64'h1260000000000000;
    #10 assign a = 64'h2D9FFFFFFFFFFFFF; assign b = 64'h126FFFFFFFFFFFFF;

    #10 $display("\n2**-293 * 2**-730:");
    #10 assign a = 64'h2DA0000000000000; assign b = 64'h1250000000000000;
    #10 assign a = 64'h2DAFFFFFFFFFFFFF; assign b = 64'h125FFFFFFFFFFFFF;

    #10 $display("\n2**-292 * 2**-731:");
    #10 assign a = 64'h2DB0000000000000; assign b = 64'h1240000000000000;
    #10 assign a = 64'h2DBFFFFFFFFFFFFF; assign b = 64'h124FFFFFFFFFFFFF;

    #10 $display("\n2**-291 * 2**-732:");
    #10 assign a = 64'h2DC0000000000000; assign b = 64'h1230000000000000;
    #10 assign a = 64'h2DCFFFFFFFFFFFFF; assign b = 64'h123FFFFFFFFFFFFF;

    #10 $display("\n2**-290 * 2**-733:");
    #10 assign a = 64'h2DD0000000000000; assign b = 64'h1220000000000000;
    #10 assign a = 64'h2DDFFFFFFFFFFFFF; assign b = 64'h122FFFFFFFFFFFFF;

    #10 $display("\n2**-289 * 2**-734:");
    #10 assign a = 64'h2DE0000000000000; assign b = 64'h1210000000000000;
    #10 assign a = 64'h2DEFFFFFFFFFFFFF; assign b = 64'h121FFFFFFFFFFFFF;

    #10 $display("\n2**-288 * 2**-735:");
    #10 assign a = 64'h2DF0000000000000; assign b = 64'h1200000000000000;
    #10 assign a = 64'h2DFFFFFFFFFFFFFF; assign b = 64'h120FFFFFFFFFFFFF;

    #10 $display("\n2**-287 * 2**-736:");
    #10 assign a = 64'h2E00000000000000; assign b = 64'h11F0000000000000;
    #10 assign a = 64'h2E0FFFFFFFFFFFFF; assign b = 64'h11FFFFFFFFFFFFFF;

    #10 $display("\n2**-286 * 2**-737:");
    #10 assign a = 64'h2E10000000000000; assign b = 64'h11E0000000000000;
    #10 assign a = 64'h2E1FFFFFFFFFFFFF; assign b = 64'h11EFFFFFFFFFFFFF;

    #10 $display("\n2**-285 * 2**-738:");
    #10 assign a = 64'h2E20000000000000; assign b = 64'h11D0000000000000;
    #10 assign a = 64'h2E2FFFFFFFFFFFFF; assign b = 64'h11DFFFFFFFFFFFFF;

    #10 $display("\n2**-284 * 2**-739:");
    #10 assign a = 64'h2E30000000000000; assign b = 64'h11C0000000000000;
    #10 assign a = 64'h2E3FFFFFFFFFFFFF; assign b = 64'h11CFFFFFFFFFFFFF;

    #10 $display("\n2**-283 * 2**-740:");
    #10 assign a = 64'h2E40000000000000; assign b = 64'h11B0000000000000;
    #10 assign a = 64'h2E4FFFFFFFFFFFFF; assign b = 64'h11BFFFFFFFFFFFFF;

    #10 $display("\n2**-282 * 2**-741:");
    #10 assign a = 64'h2E50000000000000; assign b = 64'h11A0000000000000;
    #10 assign a = 64'h2E5FFFFFFFFFFFFF; assign b = 64'h11AFFFFFFFFFFFFF;

    #10 $display("\n2**-281 * 2**-742:");
    #10 assign a = 64'h2E60000000000000; assign b = 64'h1190000000000000;
    #10 assign a = 64'h2E6FFFFFFFFFFFFF; assign b = 64'h119FFFFFFFFFFFFF;

    #10 $display("\n2**-280 * 2**-743:");
    #10 assign a = 64'h2E70000000000000; assign b = 64'h1180000000000000;
    #10 assign a = 64'h2E7FFFFFFFFFFFFF; assign b = 64'h118FFFFFFFFFFFFF;

    #10 $display("\n2**-279 * 2**-744:");
    #10 assign a = 64'h2E80000000000000; assign b = 64'h1170000000000000;
    #10 assign a = 64'h2E8FFFFFFFFFFFFF; assign b = 64'h117FFFFFFFFFFFFF;

    #10 $display("\n2**-278 * 2**-745:");
    #10 assign a = 64'h2E90000000000000; assign b = 64'h1160000000000000;
    #10 assign a = 64'h2E9FFFFFFFFFFFFF; assign b = 64'h116FFFFFFFFFFFFF;

    #10 $display("\n2**-277 * 2**-746:");
    #10 assign a = 64'h2EA0000000000000; assign b = 64'h1150000000000000;
    #10 assign a = 64'h2EAFFFFFFFFFFFFF; assign b = 64'h115FFFFFFFFFFFFF;

    #10 $display("\n2**-276 * 2**-747:");
    #10 assign a = 64'h2EB0000000000000; assign b = 64'h1140000000000000;
    #10 assign a = 64'h2EBFFFFFFFFFFFFF; assign b = 64'h114FFFFFFFFFFFFF;

    #10 $display("\n2**-275 * 2**-748:");
    #10 assign a = 64'h2EC0000000000000; assign b = 64'h1130000000000000;
    #10 assign a = 64'h2ECFFFFFFFFFFFFF; assign b = 64'h113FFFFFFFFFFFFF;

    #10 $display("\n2**-274 * 2**-749:");
    #10 assign a = 64'h2ED0000000000000; assign b = 64'h1120000000000000;
    #10 assign a = 64'h2EDFFFFFFFFFFFFF; assign b = 64'h112FFFFFFFFFFFFF;

    #10 $display("\n2**-273 * 2**-750:");
    #10 assign a = 64'h2EE0000000000000; assign b = 64'h1110000000000000;
    #10 assign a = 64'h2EEFFFFFFFFFFFFF; assign b = 64'h111FFFFFFFFFFFFF;

    #10 $display("\n2**-272 * 2**-751:");
    #10 assign a = 64'h2EF0000000000000; assign b = 64'h1100000000000000;
    #10 assign a = 64'h2EFFFFFFFFFFFFFF; assign b = 64'h110FFFFFFFFFFFFF;

    #10 $display("\n2**-271 * 2**-752:");
    #10 assign a = 64'h2F00000000000000; assign b = 64'h10F0000000000000;
    #10 assign a = 64'h2F0FFFFFFFFFFFFF; assign b = 64'h10FFFFFFFFFFFFFF;

    #10 $display("\n2**-270 * 2**-753:");
    #10 assign a = 64'h2F10000000000000; assign b = 64'h10E0000000000000;
    #10 assign a = 64'h2F1FFFFFFFFFFFFF; assign b = 64'h10EFFFFFFFFFFFFF;

    #10 $display("\n2**-269 * 2**-754:");
    #10 assign a = 64'h2F20000000000000; assign b = 64'h10D0000000000000;
    #10 assign a = 64'h2F2FFFFFFFFFFFFF; assign b = 64'h10DFFFFFFFFFFFFF;

    #10 $display("\n2**-268 * 2**-755:");
    #10 assign a = 64'h2F30000000000000; assign b = 64'h10C0000000000000;
    #10 assign a = 64'h2F3FFFFFFFFFFFFF; assign b = 64'h10CFFFFFFFFFFFFF;

    #10 $display("\n2**-267 * 2**-756:");
    #10 assign a = 64'h2F40000000000000; assign b = 64'h10B0000000000000;
    #10 assign a = 64'h2F4FFFFFFFFFFFFF; assign b = 64'h10BFFFFFFFFFFFFF;

    #10 $display("\n2**-266 * 2**-757:");
    #10 assign a = 64'h2F50000000000000; assign b = 64'h10A0000000000000;
    #10 assign a = 64'h2F5FFFFFFFFFFFFF; assign b = 64'h10AFFFFFFFFFFFFF;

    #10 $display("\n2**-265 * 2**-758:");
    #10 assign a = 64'h2F60000000000000; assign b = 64'h1090000000000000;
    #10 assign a = 64'h2F6FFFFFFFFFFFFF; assign b = 64'h109FFFFFFFFFFFFF;

    #10 $display("\n2**-264 * 2**-759:");
    #10 assign a = 64'h2F70000000000000; assign b = 64'h1080000000000000;
    #10 assign a = 64'h2F7FFFFFFFFFFFFF; assign b = 64'h108FFFFFFFFFFFFF;

    #10 $display("\n2**-263 * 2**-760:");
    #10 assign a = 64'h2F80000000000000; assign b = 64'h1070000000000000;
    #10 assign a = 64'h2F8FFFFFFFFFFFFF; assign b = 64'h107FFFFFFFFFFFFF;

    #10 $display("\n2**-262 * 2**-761:");
    #10 assign a = 64'h2F90000000000000; assign b = 64'h1060000000000000;
    #10 assign a = 64'h2F9FFFFFFFFFFFFF; assign b = 64'h106FFFFFFFFFFFFF;

    #10 $display("\n2**-261 * 2**-762:");
    #10 assign a = 64'h2FA0000000000000; assign b = 64'h1050000000000000;
    #10 assign a = 64'h2FAFFFFFFFFFFFFF; assign b = 64'h105FFFFFFFFFFFFF;

    #10 $display("\n2**-260 * 2**-763:");
    #10 assign a = 64'h2FB0000000000000; assign b = 64'h1040000000000000;
    #10 assign a = 64'h2FBFFFFFFFFFFFFF; assign b = 64'h104FFFFFFFFFFFFF;

    #10 $display("\n2**-259 * 2**-764:");
    #10 assign a = 64'h2FC0000000000000; assign b = 64'h1030000000000000;
    #10 assign a = 64'h2FCFFFFFFFFFFFFF; assign b = 64'h103FFFFFFFFFFFFF;

    #10 $display("\n2**-258 * 2**-765:");
    #10 assign a = 64'h2FD0000000000000; assign b = 64'h1020000000000000;
    #10 assign a = 64'h2FDFFFFFFFFFFFFF; assign b = 64'h102FFFFFFFFFFFFF;

    #10 $display("\n2**-257 * 2**-766:");
    #10 assign a = 64'h2FE0000000000000; assign b = 64'h1010000000000000;
    #10 assign a = 64'h2FEFFFFFFFFFFFFF; assign b = 64'h101FFFFFFFFFFFFF;

    #10 $display("\n2**-256 * 2**-767:");
    #10 assign a = 64'h2FF0000000000000; assign b = 64'h1000000000000000;
    #10 assign a = 64'h2FFFFFFFFFFFFFFF; assign b = 64'h100FFFFFFFFFFFFF;

    #10 $display("\n2**-255 * 2**-768:");
    #10 assign a = 64'h3000000000000000; assign b = 64'h0FF0000000000000;
    #10 assign a = 64'h300FFFFFFFFFFFFF; assign b = 64'h0FFFFFFFFFFFFFFF;

    #10 $display("\n2**-254 * 2**-769:");
    #10 assign a = 64'h3010000000000000; assign b = 64'h0FE0000000000000;
    #10 assign a = 64'h301FFFFFFFFFFFFF; assign b = 64'h0FEFFFFFFFFFFFFF;

    #10 $display("\n2**-253 * 2**-770:");
    #10 assign a = 64'h3020000000000000; assign b = 64'h0FD0000000000000;
    #10 assign a = 64'h302FFFFFFFFFFFFF; assign b = 64'h0FDFFFFFFFFFFFFF;

    #10 $display("\n2**-252 * 2**-771:");
    #10 assign a = 64'h3030000000000000; assign b = 64'h0FC0000000000000;
    #10 assign a = 64'h303FFFFFFFFFFFFF; assign b = 64'h0FCFFFFFFFFFFFFF;

    #10 $display("\n2**-251 * 2**-772:");
    #10 assign a = 64'h3040000000000000; assign b = 64'h0FB0000000000000;
    #10 assign a = 64'h304FFFFFFFFFFFFF; assign b = 64'h0FBFFFFFFFFFFFFF;

    #10 $display("\n2**-250 * 2**-773:");
    #10 assign a = 64'h3050000000000000; assign b = 64'h0FA0000000000000;
    #10 assign a = 64'h305FFFFFFFFFFFFF; assign b = 64'h0FAFFFFFFFFFFFFF;

    #10 $display("\n2**-249 * 2**-774:");
    #10 assign a = 64'h3060000000000000; assign b = 64'h0F90000000000000;
    #10 assign a = 64'h306FFFFFFFFFFFFF; assign b = 64'h0F9FFFFFFFFFFFFF;

    #10 $display("\n2**-248 * 2**-775:");
    #10 assign a = 64'h3070000000000000; assign b = 64'h0F80000000000000;
    #10 assign a = 64'h307FFFFFFFFFFFFF; assign b = 64'h0F8FFFFFFFFFFFFF;

    #10 $display("\n2**-247 * 2**-776:");
    #10 assign a = 64'h3080000000000000; assign b = 64'h0F70000000000000;
    #10 assign a = 64'h308FFFFFFFFFFFFF; assign b = 64'h0F7FFFFFFFFFFFFF;

    #10 $display("\n2**-246 * 2**-777:");
    #10 assign a = 64'h3090000000000000; assign b = 64'h0F60000000000000;
    #10 assign a = 64'h309FFFFFFFFFFFFF; assign b = 64'h0F6FFFFFFFFFFFFF;

    #10 $display("\n2**-245 * 2**-778:");
    #10 assign a = 64'h30A0000000000000; assign b = 64'h0F50000000000000;
    #10 assign a = 64'h30AFFFFFFFFFFFFF; assign b = 64'h0F5FFFFFFFFFFFFF;

    #10 $display("\n2**-244 * 2**-779:");
    #10 assign a = 64'h30B0000000000000; assign b = 64'h0F40000000000000;
    #10 assign a = 64'h30BFFFFFFFFFFFFF; assign b = 64'h0F4FFFFFFFFFFFFF;

    #10 $display("\n2**-243 * 2**-780:");
    #10 assign a = 64'h30C0000000000000; assign b = 64'h0F30000000000000;
    #10 assign a = 64'h30CFFFFFFFFFFFFF; assign b = 64'h0F3FFFFFFFFFFFFF;

    #10 $display("\n2**-242 * 2**-781:");
    #10 assign a = 64'h30D0000000000000; assign b = 64'h0F20000000000000;
    #10 assign a = 64'h30DFFFFFFFFFFFFF; assign b = 64'h0F2FFFFFFFFFFFFF;

    #10 $display("\n2**-241 * 2**-782:");
    #10 assign a = 64'h30E0000000000000; assign b = 64'h0F10000000000000;
    #10 assign a = 64'h30EFFFFFFFFFFFFF; assign b = 64'h0F1FFFFFFFFFFFFF;

    #10 $display("\n2**-240 * 2**-783:");
    #10 assign a = 64'h30F0000000000000; assign b = 64'h0F00000000000000;
    #10 assign a = 64'h30FFFFFFFFFFFFFF; assign b = 64'h0F0FFFFFFFFFFFFF;

    #10 $display("\n2**-239 * 2**-784:");
    #10 assign a = 64'h3100000000000000; assign b = 64'h0EF0000000000000;
    #10 assign a = 64'h310FFFFFFFFFFFFF; assign b = 64'h0EFFFFFFFFFFFFFF;

    #10 $display("\n2**-238 * 2**-785:");
    #10 assign a = 64'h3110000000000000; assign b = 64'h0EE0000000000000;
    #10 assign a = 64'h311FFFFFFFFFFFFF; assign b = 64'h0EEFFFFFFFFFFFFF;

    #10 $display("\n2**-237 * 2**-786:");
    #10 assign a = 64'h3120000000000000; assign b = 64'h0ED0000000000000;
    #10 assign a = 64'h312FFFFFFFFFFFFF; assign b = 64'h0EDFFFFFFFFFFFFF;

    #10 $display("\n2**-236 * 2**-787:");
    #10 assign a = 64'h3130000000000000; assign b = 64'h0EC0000000000000;
    #10 assign a = 64'h313FFFFFFFFFFFFF; assign b = 64'h0ECFFFFFFFFFFFFF;

    #10 $display("\n2**-235 * 2**-788:");
    #10 assign a = 64'h3140000000000000; assign b = 64'h0EB0000000000000;
    #10 assign a = 64'h314FFFFFFFFFFFFF; assign b = 64'h0EBFFFFFFFFFFFFF;

    #10 $display("\n2**-234 * 2**-789:");
    #10 assign a = 64'h3150000000000000; assign b = 64'h0EA0000000000000;
    #10 assign a = 64'h315FFFFFFFFFFFFF; assign b = 64'h0EAFFFFFFFFFFFFF;

    #10 $display("\n2**-233 * 2**-790:");
    #10 assign a = 64'h3160000000000000; assign b = 64'h0E90000000000000;
    #10 assign a = 64'h316FFFFFFFFFFFFF; assign b = 64'h0E9FFFFFFFFFFFFF;

    #10 $display("\n2**-232 * 2**-791:");
    #10 assign a = 64'h3170000000000000; assign b = 64'h0E80000000000000;
    #10 assign a = 64'h317FFFFFFFFFFFFF; assign b = 64'h0E8FFFFFFFFFFFFF;

    #10 $display("\n2**-231 * 2**-792:");
    #10 assign a = 64'h3180000000000000; assign b = 64'h0E70000000000000;
    #10 assign a = 64'h318FFFFFFFFFFFFF; assign b = 64'h0E7FFFFFFFFFFFFF;

    #10 $display("\n2**-230 * 2**-793:");
    #10 assign a = 64'h3190000000000000; assign b = 64'h0E60000000000000;
    #10 assign a = 64'h319FFFFFFFFFFFFF; assign b = 64'h0E6FFFFFFFFFFFFF;

    #10 $display("\n2**-229 * 2**-794:");
    #10 assign a = 64'h31A0000000000000; assign b = 64'h0E50000000000000;
    #10 assign a = 64'h31AFFFFFFFFFFFFF; assign b = 64'h0E5FFFFFFFFFFFFF;

    #10 $display("\n2**-228 * 2**-795:");
    #10 assign a = 64'h31B0000000000000; assign b = 64'h0E40000000000000;
    #10 assign a = 64'h31BFFFFFFFFFFFFF; assign b = 64'h0E4FFFFFFFFFFFFF;

    #10 $display("\n2**-227 * 2**-796:");
    #10 assign a = 64'h31C0000000000000; assign b = 64'h0E30000000000000;
    #10 assign a = 64'h31CFFFFFFFFFFFFF; assign b = 64'h0E3FFFFFFFFFFFFF;

    #10 $display("\n2**-226 * 2**-797:");
    #10 assign a = 64'h31D0000000000000; assign b = 64'h0E20000000000000;
    #10 assign a = 64'h31DFFFFFFFFFFFFF; assign b = 64'h0E2FFFFFFFFFFFFF;

    #10 $display("\n2**-225 * 2**-798:");
    #10 assign a = 64'h31E0000000000000; assign b = 64'h0E10000000000000;
    #10 assign a = 64'h31EFFFFFFFFFFFFF; assign b = 64'h0E1FFFFFFFFFFFFF;

    #10 $display("\n2**-224 * 2**-799:");
    #10 assign a = 64'h31F0000000000000; assign b = 64'h0E00000000000000;
    #10 assign a = 64'h31FFFFFFFFFFFFFF; assign b = 64'h0E0FFFFFFFFFFFFF;

    #10 $display("\n2**-223 * 2**-800:");
    #10 assign a = 64'h3200000000000000; assign b = 64'h0DF0000000000000;
    #10 assign a = 64'h320FFFFFFFFFFFFF; assign b = 64'h0DFFFFFFFFFFFFFF;

    #10 $display("\n2**-222 * 2**-801:");
    #10 assign a = 64'h3210000000000000; assign b = 64'h0DE0000000000000;
    #10 assign a = 64'h321FFFFFFFFFFFFF; assign b = 64'h0DEFFFFFFFFFFFFF;

    #10 $display("\n2**-221 * 2**-802:");
    #10 assign a = 64'h3220000000000000; assign b = 64'h0DD0000000000000;
    #10 assign a = 64'h322FFFFFFFFFFFFF; assign b = 64'h0DDFFFFFFFFFFFFF;

    #10 $display("\n2**-220 * 2**-803:");
    #10 assign a = 64'h3230000000000000; assign b = 64'h0DC0000000000000;
    #10 assign a = 64'h323FFFFFFFFFFFFF; assign b = 64'h0DCFFFFFFFFFFFFF;

    #10 $display("\n2**-219 * 2**-804:");
    #10 assign a = 64'h3240000000000000; assign b = 64'h0DB0000000000000;
    #10 assign a = 64'h324FFFFFFFFFFFFF; assign b = 64'h0DBFFFFFFFFFFFFF;

    #10 $display("\n2**-218 * 2**-805:");
    #10 assign a = 64'h3250000000000000; assign b = 64'h0DA0000000000000;
    #10 assign a = 64'h325FFFFFFFFFFFFF; assign b = 64'h0DAFFFFFFFFFFFFF;

    #10 $display("\n2**-217 * 2**-806:");
    #10 assign a = 64'h3260000000000000; assign b = 64'h0D90000000000000;
    #10 assign a = 64'h326FFFFFFFFFFFFF; assign b = 64'h0D9FFFFFFFFFFFFF;

    #10 $display("\n2**-216 * 2**-807:");
    #10 assign a = 64'h3270000000000000; assign b = 64'h0D80000000000000;
    #10 assign a = 64'h327FFFFFFFFFFFFF; assign b = 64'h0D8FFFFFFFFFFFFF;

    #10 $display("\n2**-215 * 2**-808:");
    #10 assign a = 64'h3280000000000000; assign b = 64'h0D70000000000000;
    #10 assign a = 64'h328FFFFFFFFFFFFF; assign b = 64'h0D7FFFFFFFFFFFFF;

    #10 $display("\n2**-214 * 2**-809:");
    #10 assign a = 64'h3290000000000000; assign b = 64'h0D60000000000000;
    #10 assign a = 64'h329FFFFFFFFFFFFF; assign b = 64'h0D6FFFFFFFFFFFFF;

    #10 $display("\n2**-213 * 2**-810:");
    #10 assign a = 64'h32A0000000000000; assign b = 64'h0D50000000000000;
    #10 assign a = 64'h32AFFFFFFFFFFFFF; assign b = 64'h0D5FFFFFFFFFFFFF;

    #10 $display("\n2**-212 * 2**-811:");
    #10 assign a = 64'h32B0000000000000; assign b = 64'h0D40000000000000;
    #10 assign a = 64'h32BFFFFFFFFFFFFF; assign b = 64'h0D4FFFFFFFFFFFFF;

    #10 $display("\n2**-211 * 2**-812:");
    #10 assign a = 64'h32C0000000000000; assign b = 64'h0D30000000000000;
    #10 assign a = 64'h32CFFFFFFFFFFFFF; assign b = 64'h0D3FFFFFFFFFFFFF;

    #10 $display("\n2**-210 * 2**-813:");
    #10 assign a = 64'h32D0000000000000; assign b = 64'h0D20000000000000;
    #10 assign a = 64'h32DFFFFFFFFFFFFF; assign b = 64'h0D2FFFFFFFFFFFFF;

    #10 $display("\n2**-209 * 2**-814:");
    #10 assign a = 64'h32E0000000000000; assign b = 64'h0D10000000000000;
    #10 assign a = 64'h32EFFFFFFFFFFFFF; assign b = 64'h0D1FFFFFFFFFFFFF;

    #10 $display("\n2**-208 * 2**-815:");
    #10 assign a = 64'h32F0000000000000; assign b = 64'h0D00000000000000;
    #10 assign a = 64'h32FFFFFFFFFFFFFF; assign b = 64'h0D0FFFFFFFFFFFFF;

    #10 $display("\n2**-207 * 2**-816:");
    #10 assign a = 64'h3300000000000000; assign b = 64'h0CF0000000000000;
    #10 assign a = 64'h330FFFFFFFFFFFFF; assign b = 64'h0CFFFFFFFFFFFFFF;

    #10 $display("\n2**-206 * 2**-817:");
    #10 assign a = 64'h3310000000000000; assign b = 64'h0CE0000000000000;
    #10 assign a = 64'h331FFFFFFFFFFFFF; assign b = 64'h0CEFFFFFFFFFFFFF;

    #10 $display("\n2**-205 * 2**-818:");
    #10 assign a = 64'h3320000000000000; assign b = 64'h0CD0000000000000;
    #10 assign a = 64'h332FFFFFFFFFFFFF; assign b = 64'h0CDFFFFFFFFFFFFF;

    #10 $display("\n2**-204 * 2**-819:");
    #10 assign a = 64'h3330000000000000; assign b = 64'h0CC0000000000000;
    #10 assign a = 64'h333FFFFFFFFFFFFF; assign b = 64'h0CCFFFFFFFFFFFFF;

    #10 $display("\n2**-203 * 2**-820:");
    #10 assign a = 64'h3340000000000000; assign b = 64'h0CB0000000000000;
    #10 assign a = 64'h334FFFFFFFFFFFFF; assign b = 64'h0CBFFFFFFFFFFFFF;

    #10 $display("\n2**-202 * 2**-821:");
    #10 assign a = 64'h3350000000000000; assign b = 64'h0CA0000000000000;
    #10 assign a = 64'h335FFFFFFFFFFFFF; assign b = 64'h0CAFFFFFFFFFFFFF;

    #10 $display("\n2**-201 * 2**-822:");
    #10 assign a = 64'h3360000000000000; assign b = 64'h0C90000000000000;
    #10 assign a = 64'h336FFFFFFFFFFFFF; assign b = 64'h0C9FFFFFFFFFFFFF;

    #10 $display("\n2**-200 * 2**-823:");
    #10 assign a = 64'h3370000000000000; assign b = 64'h0C80000000000000;
    #10 assign a = 64'h337FFFFFFFFFFFFF; assign b = 64'h0C8FFFFFFFFFFFFF;

    #10 $display("\n2**-199 * 2**-824:");
    #10 assign a = 64'h3380000000000000; assign b = 64'h0C70000000000000;
    #10 assign a = 64'h338FFFFFFFFFFFFF; assign b = 64'h0C7FFFFFFFFFFFFF;

    #10 $display("\n2**-198 * 2**-825:");
    #10 assign a = 64'h3390000000000000; assign b = 64'h0C60000000000000;
    #10 assign a = 64'h339FFFFFFFFFFFFF; assign b = 64'h0C6FFFFFFFFFFFFF;

    #10 $display("\n2**-197 * 2**-826:");
    #10 assign a = 64'h33A0000000000000; assign b = 64'h0C50000000000000;
    #10 assign a = 64'h33AFFFFFFFFFFFFF; assign b = 64'h0C5FFFFFFFFFFFFF;

    #10 $display("\n2**-196 * 2**-827:");
    #10 assign a = 64'h33B0000000000000; assign b = 64'h0C40000000000000;
    #10 assign a = 64'h33BFFFFFFFFFFFFF; assign b = 64'h0C4FFFFFFFFFFFFF;

    #10 $display("\n2**-195 * 2**-828:");
    #10 assign a = 64'h33C0000000000000; assign b = 64'h0C30000000000000;
    #10 assign a = 64'h33CFFFFFFFFFFFFF; assign b = 64'h0C3FFFFFFFFFFFFF;

    #10 $display("\n2**-194 * 2**-829:");
    #10 assign a = 64'h33D0000000000000; assign b = 64'h0C20000000000000;
    #10 assign a = 64'h33DFFFFFFFFFFFFF; assign b = 64'h0C2FFFFFFFFFFFFF;

    #10 $display("\n2**-193 * 2**-830:");
    #10 assign a = 64'h33E0000000000000; assign b = 64'h0C10000000000000;
    #10 assign a = 64'h33EFFFFFFFFFFFFF; assign b = 64'h0C1FFFFFFFFFFFFF;

    #10 $display("\n2**-192 * 2**-831:");
    #10 assign a = 64'h33F0000000000000; assign b = 64'h0C00000000000000;
    #10 assign a = 64'h33FFFFFFFFFFFFFF; assign b = 64'h0C0FFFFFFFFFFFFF;

    #10 $display("\n2**-191 * 2**-832:");
    #10 assign a = 64'h3400000000000000; assign b = 64'h0BF0000000000000;
    #10 assign a = 64'h340FFFFFFFFFFFFF; assign b = 64'h0BFFFFFFFFFFFFFF;

    #10 $display("\n2**-190 * 2**-833:");
    #10 assign a = 64'h3410000000000000; assign b = 64'h0BE0000000000000;
    #10 assign a = 64'h341FFFFFFFFFFFFF; assign b = 64'h0BEFFFFFFFFFFFFF;

    #10 $display("\n2**-189 * 2**-834:");
    #10 assign a = 64'h3420000000000000; assign b = 64'h0BD0000000000000;
    #10 assign a = 64'h342FFFFFFFFFFFFF; assign b = 64'h0BDFFFFFFFFFFFFF;

    #10 $display("\n2**-188 * 2**-835:");
    #10 assign a = 64'h3430000000000000; assign b = 64'h0BC0000000000000;
    #10 assign a = 64'h343FFFFFFFFFFFFF; assign b = 64'h0BCFFFFFFFFFFFFF;

    #10 $display("\n2**-187 * 2**-836:");
    #10 assign a = 64'h3440000000000000; assign b = 64'h0BB0000000000000;
    #10 assign a = 64'h344FFFFFFFFFFFFF; assign b = 64'h0BBFFFFFFFFFFFFF;

    #10 $display("\n2**-186 * 2**-837:");
    #10 assign a = 64'h3450000000000000; assign b = 64'h0BA0000000000000;
    #10 assign a = 64'h345FFFFFFFFFFFFF; assign b = 64'h0BAFFFFFFFFFFFFF;

    #10 $display("\n2**-185 * 2**-838:");
    #10 assign a = 64'h3460000000000000; assign b = 64'h0B90000000000000;
    #10 assign a = 64'h346FFFFFFFFFFFFF; assign b = 64'h0B9FFFFFFFFFFFFF;

    #10 $display("\n2**-184 * 2**-839:");
    #10 assign a = 64'h3470000000000000; assign b = 64'h0B80000000000000;
    #10 assign a = 64'h347FFFFFFFFFFFFF; assign b = 64'h0B8FFFFFFFFFFFFF;

    #10 $display("\n2**-183 * 2**-840:");
    #10 assign a = 64'h3480000000000000; assign b = 64'h0B70000000000000;
    #10 assign a = 64'h348FFFFFFFFFFFFF; assign b = 64'h0B7FFFFFFFFFFFFF;

    #10 $display("\n2**-182 * 2**-841:");
    #10 assign a = 64'h3490000000000000; assign b = 64'h0B60000000000000;
    #10 assign a = 64'h349FFFFFFFFFFFFF; assign b = 64'h0B6FFFFFFFFFFFFF;

    #10 $display("\n2**-181 * 2**-842:");
    #10 assign a = 64'h34A0000000000000; assign b = 64'h0B50000000000000;
    #10 assign a = 64'h34AFFFFFFFFFFFFF; assign b = 64'h0B5FFFFFFFFFFFFF;

    #10 $display("\n2**-180 * 2**-843:");
    #10 assign a = 64'h34B0000000000000; assign b = 64'h0B40000000000000;
    #10 assign a = 64'h34BFFFFFFFFFFFFF; assign b = 64'h0B4FFFFFFFFFFFFF;

    #10 $display("\n2**-179 * 2**-844:");
    #10 assign a = 64'h34C0000000000000; assign b = 64'h0B30000000000000;
    #10 assign a = 64'h34CFFFFFFFFFFFFF; assign b = 64'h0B3FFFFFFFFFFFFF;

    #10 $display("\n2**-178 * 2**-845:");
    #10 assign a = 64'h34D0000000000000; assign b = 64'h0B20000000000000;
    #10 assign a = 64'h34DFFFFFFFFFFFFF; assign b = 64'h0B2FFFFFFFFFFFFF;

    #10 $display("\n2**-177 * 2**-846:");
    #10 assign a = 64'h34E0000000000000; assign b = 64'h0B10000000000000;
    #10 assign a = 64'h34EFFFFFFFFFFFFF; assign b = 64'h0B1FFFFFFFFFFFFF;

    #10 $display("\n2**-176 * 2**-847:");
    #10 assign a = 64'h34F0000000000000; assign b = 64'h0B00000000000000;
    #10 assign a = 64'h34FFFFFFFFFFFFFF; assign b = 64'h0B0FFFFFFFFFFFFF;

    #10 $display("\n2**-175 * 2**-848:");
    #10 assign a = 64'h3500000000000000; assign b = 64'h0AF0000000000000;
    #10 assign a = 64'h350FFFFFFFFFFFFF; assign b = 64'h0AFFFFFFFFFFFFFF;

    #10 $display("\n2**-174 * 2**-849:");
    #10 assign a = 64'h3510000000000000; assign b = 64'h0AE0000000000000;
    #10 assign a = 64'h351FFFFFFFFFFFFF; assign b = 64'h0AEFFFFFFFFFFFFF;

    #10 $display("\n2**-173 * 2**-850:");
    #10 assign a = 64'h3520000000000000; assign b = 64'h0AD0000000000000;
    #10 assign a = 64'h352FFFFFFFFFFFFF; assign b = 64'h0ADFFFFFFFFFFFFF;

    #10 $display("\n2**-172 * 2**-851:");
    #10 assign a = 64'h3530000000000000; assign b = 64'h0AC0000000000000;
    #10 assign a = 64'h353FFFFFFFFFFFFF; assign b = 64'h0ACFFFFFFFFFFFFF;

    #10 $display("\n2**-171 * 2**-852:");
    #10 assign a = 64'h3540000000000000; assign b = 64'h0AB0000000000000;
    #10 assign a = 64'h354FFFFFFFFFFFFF; assign b = 64'h0ABFFFFFFFFFFFFF;

    #10 $display("\n2**-170 * 2**-853:");
    #10 assign a = 64'h3550000000000000; assign b = 64'h0AA0000000000000;
    #10 assign a = 64'h355FFFFFFFFFFFFF; assign b = 64'h0AAFFFFFFFFFFFFF;

    #10 $display("\n2**-169 * 2**-854:");
    #10 assign a = 64'h3560000000000000; assign b = 64'h0A90000000000000;
    #10 assign a = 64'h356FFFFFFFFFFFFF; assign b = 64'h0A9FFFFFFFFFFFFF;

    #10 $display("\n2**-168 * 2**-855:");
    #10 assign a = 64'h3570000000000000; assign b = 64'h0A80000000000000;
    #10 assign a = 64'h357FFFFFFFFFFFFF; assign b = 64'h0A8FFFFFFFFFFFFF;

    #10 $display("\n2**-167 * 2**-856:");
    #10 assign a = 64'h3580000000000000; assign b = 64'h0A70000000000000;
    #10 assign a = 64'h358FFFFFFFFFFFFF; assign b = 64'h0A7FFFFFFFFFFFFF;

    #10 $display("\n2**-166 * 2**-857:");
    #10 assign a = 64'h3590000000000000; assign b = 64'h0A60000000000000;
    #10 assign a = 64'h359FFFFFFFFFFFFF; assign b = 64'h0A6FFFFFFFFFFFFF;

    #10 $display("\n2**-165 * 2**-858:");
    #10 assign a = 64'h35A0000000000000; assign b = 64'h0A50000000000000;
    #10 assign a = 64'h35AFFFFFFFFFFFFF; assign b = 64'h0A5FFFFFFFFFFFFF;

    #10 $display("\n2**-164 * 2**-859:");
    #10 assign a = 64'h35B0000000000000; assign b = 64'h0A40000000000000;
    #10 assign a = 64'h35BFFFFFFFFFFFFF; assign b = 64'h0A4FFFFFFFFFFFFF;

    #10 $display("\n2**-163 * 2**-860:");
    #10 assign a = 64'h35C0000000000000; assign b = 64'h0A30000000000000;
    #10 assign a = 64'h35CFFFFFFFFFFFFF; assign b = 64'h0A3FFFFFFFFFFFFF;

    #10 $display("\n2**-162 * 2**-861:");
    #10 assign a = 64'h35D0000000000000; assign b = 64'h0A20000000000000;
    #10 assign a = 64'h35DFFFFFFFFFFFFF; assign b = 64'h0A2FFFFFFFFFFFFF;

    #10 $display("\n2**-161 * 2**-862:");
    #10 assign a = 64'h35E0000000000000; assign b = 64'h0A10000000000000;
    #10 assign a = 64'h35EFFFFFFFFFFFFF; assign b = 64'h0A1FFFFFFFFFFFFF;

    #10 $display("\n2**-160 * 2**-863:");
    #10 assign a = 64'h35F0000000000000; assign b = 64'h0A00000000000000;
    #10 assign a = 64'h35FFFFFFFFFFFFFF; assign b = 64'h0A0FFFFFFFFFFFFF;

    #10 $display("\n2**-159 * 2**-864:");
    #10 assign a = 64'h3600000000000000; assign b = 64'h09F0000000000000;
    #10 assign a = 64'h360FFFFFFFFFFFFF; assign b = 64'h09FFFFFFFFFFFFFF;

    #10 $display("\n2**-158 * 2**-865:");
    #10 assign a = 64'h3610000000000000; assign b = 64'h09E0000000000000;
    #10 assign a = 64'h361FFFFFFFFFFFFF; assign b = 64'h09EFFFFFFFFFFFFF;

    #10 $display("\n2**-157 * 2**-866:");
    #10 assign a = 64'h3620000000000000; assign b = 64'h09D0000000000000;
    #10 assign a = 64'h362FFFFFFFFFFFFF; assign b = 64'h09DFFFFFFFFFFFFF;

    #10 $display("\n2**-156 * 2**-867:");
    #10 assign a = 64'h3630000000000000; assign b = 64'h09C0000000000000;
    #10 assign a = 64'h363FFFFFFFFFFFFF; assign b = 64'h09CFFFFFFFFFFFFF;

    #10 $display("\n2**-155 * 2**-868:");
    #10 assign a = 64'h3640000000000000; assign b = 64'h09B0000000000000;
    #10 assign a = 64'h364FFFFFFFFFFFFF; assign b = 64'h09BFFFFFFFFFFFFF;

    #10 $display("\n2**-154 * 2**-869:");
    #10 assign a = 64'h3650000000000000; assign b = 64'h09A0000000000000;
    #10 assign a = 64'h365FFFFFFFFFFFFF; assign b = 64'h09AFFFFFFFFFFFFF;

    #10 $display("\n2**-153 * 2**-870:");
    #10 assign a = 64'h3660000000000000; assign b = 64'h0990000000000000;
    #10 assign a = 64'h366FFFFFFFFFFFFF; assign b = 64'h099FFFFFFFFFFFFF;

    #10 $display("\n2**-152 * 2**-871:");
    #10 assign a = 64'h3670000000000000; assign b = 64'h0980000000000000;
    #10 assign a = 64'h367FFFFFFFFFFFFF; assign b = 64'h098FFFFFFFFFFFFF;

    #10 $display("\n2**-151 * 2**-872:");
    #10 assign a = 64'h3680000000000000; assign b = 64'h0970000000000000;
    #10 assign a = 64'h368FFFFFFFFFFFFF; assign b = 64'h097FFFFFFFFFFFFF;

    #10 $display("\n2**-150 * 2**-873:");
    #10 assign a = 64'h3690000000000000; assign b = 64'h0960000000000000;
    #10 assign a = 64'h369FFFFFFFFFFFFF; assign b = 64'h096FFFFFFFFFFFFF;

    #10 $display("\n2**-149 * 2**-874:");
    #10 assign a = 64'h36A0000000000000; assign b = 64'h0950000000000000;
    #10 assign a = 64'h36AFFFFFFFFFFFFF; assign b = 64'h095FFFFFFFFFFFFF;

    #10 $display("\n2**-148 * 2**-875:");
    #10 assign a = 64'h36B0000000000000; assign b = 64'h0940000000000000;
    #10 assign a = 64'h36BFFFFFFFFFFFFF; assign b = 64'h094FFFFFFFFFFFFF;

    #10 $display("\n2**-147 * 2**-876:");
    #10 assign a = 64'h36C0000000000000; assign b = 64'h0930000000000000;
    #10 assign a = 64'h36CFFFFFFFFFFFFF; assign b = 64'h093FFFFFFFFFFFFF;

    #10 $display("\n2**-146 * 2**-877:");
    #10 assign a = 64'h36D0000000000000; assign b = 64'h0920000000000000;
    #10 assign a = 64'h36DFFFFFFFFFFFFF; assign b = 64'h092FFFFFFFFFFFFF;

    #10 $display("\n2**-145 * 2**-878:");
    #10 assign a = 64'h36E0000000000000; assign b = 64'h0910000000000000;
    #10 assign a = 64'h36EFFFFFFFFFFFFF; assign b = 64'h091FFFFFFFFFFFFF;

    #10 $display("\n2**-144 * 2**-879:");
    #10 assign a = 64'h36F0000000000000; assign b = 64'h0900000000000000;
    #10 assign a = 64'h36FFFFFFFFFFFFFF; assign b = 64'h090FFFFFFFFFFFFF;

    #10 $display("\n2**-143 * 2**-880:");
    #10 assign a = 64'h3700000000000000; assign b = 64'h08F0000000000000;
    #10 assign a = 64'h370FFFFFFFFFFFFF; assign b = 64'h08FFFFFFFFFFFFFF;

    #10 $display("\n2**-142 * 2**-881:");
    #10 assign a = 64'h3710000000000000; assign b = 64'h08E0000000000000;
    #10 assign a = 64'h371FFFFFFFFFFFFF; assign b = 64'h08EFFFFFFFFFFFFF;

    #10 $display("\n2**-141 * 2**-882:");
    #10 assign a = 64'h3720000000000000; assign b = 64'h08D0000000000000;
    #10 assign a = 64'h372FFFFFFFFFFFFF; assign b = 64'h08DFFFFFFFFFFFFF;

    #10 $display("\n2**-140 * 2**-883:");
    #10 assign a = 64'h3730000000000000; assign b = 64'h08C0000000000000;
    #10 assign a = 64'h373FFFFFFFFFFFFF; assign b = 64'h08CFFFFFFFFFFFFF;

    #10 $display("\n2**-139 * 2**-884:");
    #10 assign a = 64'h3740000000000000; assign b = 64'h08B0000000000000;
    #10 assign a = 64'h374FFFFFFFFFFFFF; assign b = 64'h08BFFFFFFFFFFFFF;

    #10 $display("\n2**-138 * 2**-885:");
    #10 assign a = 64'h3750000000000000; assign b = 64'h08A0000000000000;
    #10 assign a = 64'h375FFFFFFFFFFFFF; assign b = 64'h08AFFFFFFFFFFFFF;

    #10 $display("\n2**-137 * 2**-886:");
    #10 assign a = 64'h3760000000000000; assign b = 64'h0890000000000000;
    #10 assign a = 64'h376FFFFFFFFFFFFF; assign b = 64'h089FFFFFFFFFFFFF;

    #10 $display("\n2**-136 * 2**-887:");
    #10 assign a = 64'h3770000000000000; assign b = 64'h0880000000000000;
    #10 assign a = 64'h377FFFFFFFFFFFFF; assign b = 64'h088FFFFFFFFFFFFF;

    #10 $display("\n2**-135 * 2**-888:");
    #10 assign a = 64'h3780000000000000; assign b = 64'h0870000000000000;
    #10 assign a = 64'h378FFFFFFFFFFFFF; assign b = 64'h087FFFFFFFFFFFFF;

    #10 $display("\n2**-134 * 2**-889:");
    #10 assign a = 64'h3790000000000000; assign b = 64'h0860000000000000;
    #10 assign a = 64'h379FFFFFFFFFFFFF; assign b = 64'h086FFFFFFFFFFFFF;

    #10 $display("\n2**-133 * 2**-890:");
    #10 assign a = 64'h37A0000000000000; assign b = 64'h0850000000000000;
    #10 assign a = 64'h37AFFFFFFFFFFFFF; assign b = 64'h085FFFFFFFFFFFFF;

    #10 $display("\n2**-132 * 2**-891:");
    #10 assign a = 64'h37B0000000000000; assign b = 64'h0840000000000000;
    #10 assign a = 64'h37BFFFFFFFFFFFFF; assign b = 64'h084FFFFFFFFFFFFF;

    #10 $display("\n2**-131 * 2**-892:");
    #10 assign a = 64'h37C0000000000000; assign b = 64'h0830000000000000;
    #10 assign a = 64'h37CFFFFFFFFFFFFF; assign b = 64'h083FFFFFFFFFFFFF;

    #10 $display("\n2**-130 * 2**-893:");
    #10 assign a = 64'h37D0000000000000; assign b = 64'h0820000000000000;
    #10 assign a = 64'h37DFFFFFFFFFFFFF; assign b = 64'h082FFFFFFFFFFFFF;

    #10 $display("\n2**-129 * 2**-894:");
    #10 assign a = 64'h37E0000000000000; assign b = 64'h0810000000000000;
    #10 assign a = 64'h37EFFFFFFFFFFFFF; assign b = 64'h081FFFFFFFFFFFFF;

    #10 $display("\n2**-128 * 2**-895:");
    #10 assign a = 64'h37F0000000000000; assign b = 64'h0800000000000000;
    #10 assign a = 64'h37FFFFFFFFFFFFFF; assign b = 64'h080FFFFFFFFFFFFF;

    #10 $display("\n2**-127 * 2**-896:");
    #10 assign a = 64'h3800000000000000; assign b = 64'h07F0000000000000;
    #10 assign a = 64'h380FFFFFFFFFFFFF; assign b = 64'h07FFFFFFFFFFFFFF;

    #10 $display("\n2**-126 * 2**-897:");
    #10 assign a = 64'h3810000000000000; assign b = 64'h07E0000000000000;
    #10 assign a = 64'h381FFFFFFFFFFFFF; assign b = 64'h07EFFFFFFFFFFFFF;

    #10 $display("\n2**-125 * 2**-898:");
    #10 assign a = 64'h3820000000000000; assign b = 64'h07D0000000000000;
    #10 assign a = 64'h382FFFFFFFFFFFFF; assign b = 64'h07DFFFFFFFFFFFFF;

    #10 $display("\n2**-124 * 2**-899:");
    #10 assign a = 64'h3830000000000000; assign b = 64'h07C0000000000000;
    #10 assign a = 64'h383FFFFFFFFFFFFF; assign b = 64'h07CFFFFFFFFFFFFF;

    #10 $display("\n2**-123 * 2**-900:");
    #10 assign a = 64'h3840000000000000; assign b = 64'h07B0000000000000;
    #10 assign a = 64'h384FFFFFFFFFFFFF; assign b = 64'h07BFFFFFFFFFFFFF;

    #10 $display("\n2**-122 * 2**-901:");
    #10 assign a = 64'h3850000000000000; assign b = 64'h07A0000000000000;
    #10 assign a = 64'h385FFFFFFFFFFFFF; assign b = 64'h07AFFFFFFFFFFFFF;

    #10 $display("\n2**-121 * 2**-902:");
    #10 assign a = 64'h3860000000000000; assign b = 64'h0790000000000000;
    #10 assign a = 64'h386FFFFFFFFFFFFF; assign b = 64'h079FFFFFFFFFFFFF;

    #10 $display("\n2**-120 * 2**-903:");
    #10 assign a = 64'h3870000000000000; assign b = 64'h0780000000000000;
    #10 assign a = 64'h387FFFFFFFFFFFFF; assign b = 64'h078FFFFFFFFFFFFF;

    #10 $display("\n2**-119 * 2**-904:");
    #10 assign a = 64'h3880000000000000; assign b = 64'h0770000000000000;
    #10 assign a = 64'h388FFFFFFFFFFFFF; assign b = 64'h077FFFFFFFFFFFFF;

    #10 $display("\n2**-118 * 2**-905:");
    #10 assign a = 64'h3890000000000000; assign b = 64'h0760000000000000;
    #10 assign a = 64'h389FFFFFFFFFFFFF; assign b = 64'h076FFFFFFFFFFFFF;

    #10 $display("\n2**-117 * 2**-906:");
    #10 assign a = 64'h38A0000000000000; assign b = 64'h0750000000000000;
    #10 assign a = 64'h38AFFFFFFFFFFFFF; assign b = 64'h075FFFFFFFFFFFFF;

    #10 $display("\n2**-116 * 2**-907:");
    #10 assign a = 64'h38B0000000000000; assign b = 64'h0740000000000000;
    #10 assign a = 64'h38BFFFFFFFFFFFFF; assign b = 64'h074FFFFFFFFFFFFF;

    #10 $display("\n2**-115 * 2**-908:");
    #10 assign a = 64'h38C0000000000000; assign b = 64'h0730000000000000;
    #10 assign a = 64'h38CFFFFFFFFFFFFF; assign b = 64'h073FFFFFFFFFFFFF;

    #10 $display("\n2**-114 * 2**-909:");
    #10 assign a = 64'h38D0000000000000; assign b = 64'h0720000000000000;
    #10 assign a = 64'h38DFFFFFFFFFFFFF; assign b = 64'h072FFFFFFFFFFFFF;

    #10 $display("\n2**-113 * 2**-910:");
    #10 assign a = 64'h38E0000000000000; assign b = 64'h0710000000000000;
    #10 assign a = 64'h38EFFFFFFFFFFFFF; assign b = 64'h071FFFFFFFFFFFFF;

    #10 $display("\n2**-112 * 2**-911:");
    #10 assign a = 64'h38F0000000000000; assign b = 64'h0700000000000000;
    #10 assign a = 64'h38FFFFFFFFFFFFFF; assign b = 64'h070FFFFFFFFFFFFF;

    #10 $display("\n2**-111 * 2**-912:");
    #10 assign a = 64'h3900000000000000; assign b = 64'h06F0000000000000;
    #10 assign a = 64'h390FFFFFFFFFFFFF; assign b = 64'h06FFFFFFFFFFFFFF;

    #10 $display("\n2**-110 * 2**-913:");
    #10 assign a = 64'h3910000000000000; assign b = 64'h06E0000000000000;
    #10 assign a = 64'h391FFFFFFFFFFFFF; assign b = 64'h06EFFFFFFFFFFFFF;

    #10 $display("\n2**-109 * 2**-914:");
    #10 assign a = 64'h3920000000000000; assign b = 64'h06D0000000000000;
    #10 assign a = 64'h392FFFFFFFFFFFFF; assign b = 64'h06DFFFFFFFFFFFFF;

    #10 $display("\n2**-108 * 2**-915:");
    #10 assign a = 64'h3930000000000000; assign b = 64'h06C0000000000000;
    #10 assign a = 64'h393FFFFFFFFFFFFF; assign b = 64'h06CFFFFFFFFFFFFF;

    #10 $display("\n2**-107 * 2**-916:");
    #10 assign a = 64'h3940000000000000; assign b = 64'h06B0000000000000;
    #10 assign a = 64'h394FFFFFFFFFFFFF; assign b = 64'h06BFFFFFFFFFFFFF;

    #10 $display("\n2**-106 * 2**-917:");
    #10 assign a = 64'h3950000000000000; assign b = 64'h06A0000000000000;
    #10 assign a = 64'h395FFFFFFFFFFFFF; assign b = 64'h06AFFFFFFFFFFFFF;

    #10 $display("\n2**-105 * 2**-918:");
    #10 assign a = 64'h3960000000000000; assign b = 64'h0690000000000000;
    #10 assign a = 64'h396FFFFFFFFFFFFF; assign b = 64'h069FFFFFFFFFFFFF;

    #10 $display("\n2**-104 * 2**-919:");
    #10 assign a = 64'h3970000000000000; assign b = 64'h0680000000000000;
    #10 assign a = 64'h397FFFFFFFFFFFFF; assign b = 64'h068FFFFFFFFFFFFF;

    #10 $display("\n2**-103 * 2**-920:");
    #10 assign a = 64'h3980000000000000; assign b = 64'h0670000000000000;
    #10 assign a = 64'h398FFFFFFFFFFFFF; assign b = 64'h067FFFFFFFFFFFFF;

    #10 $display("\n2**-102 * 2**-921:");
    #10 assign a = 64'h3990000000000000; assign b = 64'h0660000000000000;
    #10 assign a = 64'h399FFFFFFFFFFFFF; assign b = 64'h066FFFFFFFFFFFFF;

    #10 $display("\n2**-101 * 2**-922:");
    #10 assign a = 64'h39A0000000000000; assign b = 64'h0650000000000000;
    #10 assign a = 64'h39AFFFFFFFFFFFFF; assign b = 64'h065FFFFFFFFFFFFF;

    #10 $display("\n2**-100 * 2**-923:");
    #10 assign a = 64'h39B0000000000000; assign b = 64'h0640000000000000;
    #10 assign a = 64'h39BFFFFFFFFFFFFF; assign b = 64'h064FFFFFFFFFFFFF;

    #10 $display("\n2**-99 * 2**-924:");
    #10 assign a = 64'h39C0000000000000; assign b = 64'h0630000000000000;
    #10 assign a = 64'h39CFFFFFFFFFFFFF; assign b = 64'h063FFFFFFFFFFFFF;

    #10 $display("\n2**-98 * 2**-925:");
    #10 assign a = 64'h39D0000000000000; assign b = 64'h0620000000000000;
    #10 assign a = 64'h39DFFFFFFFFFFFFF; assign b = 64'h062FFFFFFFFFFFFF;

    #10 $display("\n2**-97 * 2**-926:");
    #10 assign a = 64'h39E0000000000000; assign b = 64'h0610000000000000;
    #10 assign a = 64'h39EFFFFFFFFFFFFF; assign b = 64'h061FFFFFFFFFFFFF;

    #10 $display("\n2**-96 * 2**-927:");
    #10 assign a = 64'h39F0000000000000; assign b = 64'h0600000000000000;
    #10 assign a = 64'h39FFFFFFFFFFFFFF; assign b = 64'h060FFFFFFFFFFFFF;

    #10 $display("\n2**-95 * 2**-928:");
    #10 assign a = 64'h3A00000000000000; assign b = 64'h05F0000000000000;
    #10 assign a = 64'h3A0FFFFFFFFFFFFF; assign b = 64'h05FFFFFFFFFFFFFF;

    #10 $display("\n2**-94 * 2**-929:");
    #10 assign a = 64'h3A10000000000000; assign b = 64'h05E0000000000000;
    #10 assign a = 64'h3A1FFFFFFFFFFFFF; assign b = 64'h05EFFFFFFFFFFFFF;

    #10 $display("\n2**-93 * 2**-930:");
    #10 assign a = 64'h3A20000000000000; assign b = 64'h05D0000000000000;
    #10 assign a = 64'h3A2FFFFFFFFFFFFF; assign b = 64'h05DFFFFFFFFFFFFF;

    #10 $display("\n2**-92 * 2**-931:");
    #10 assign a = 64'h3A30000000000000; assign b = 64'h05C0000000000000;
    #10 assign a = 64'h3A3FFFFFFFFFFFFF; assign b = 64'h05CFFFFFFFFFFFFF;

    #10 $display("\n2**-91 * 2**-932:");
    #10 assign a = 64'h3A40000000000000; assign b = 64'h05B0000000000000;
    #10 assign a = 64'h3A4FFFFFFFFFFFFF; assign b = 64'h05BFFFFFFFFFFFFF;

    #10 $display("\n2**-90 * 2**-933:");
    #10 assign a = 64'h3A50000000000000; assign b = 64'h05A0000000000000;
    #10 assign a = 64'h3A5FFFFFFFFFFFFF; assign b = 64'h05AFFFFFFFFFFFFF;

    #10 $display("\n2**-89 * 2**-934:");
    #10 assign a = 64'h3A60000000000000; assign b = 64'h0590000000000000;
    #10 assign a = 64'h3A6FFFFFFFFFFFFF; assign b = 64'h059FFFFFFFFFFFFF;

    #10 $display("\n2**-88 * 2**-935:");
    #10 assign a = 64'h3A70000000000000; assign b = 64'h0580000000000000;
    #10 assign a = 64'h3A7FFFFFFFFFFFFF; assign b = 64'h058FFFFFFFFFFFFF;

    #10 $display("\n2**-87 * 2**-936:");
    #10 assign a = 64'h3A80000000000000; assign b = 64'h0570000000000000;
    #10 assign a = 64'h3A8FFFFFFFFFFFFF; assign b = 64'h057FFFFFFFFFFFFF;

    #10 $display("\n2**-86 * 2**-937:");
    #10 assign a = 64'h3A90000000000000; assign b = 64'h0560000000000000;
    #10 assign a = 64'h3A9FFFFFFFFFFFFF; assign b = 64'h056FFFFFFFFFFFFF;

    #10 $display("\n2**-85 * 2**-938:");
    #10 assign a = 64'h3AA0000000000000; assign b = 64'h0550000000000000;
    #10 assign a = 64'h3AAFFFFFFFFFFFFF; assign b = 64'h055FFFFFFFFFFFFF;

    #10 $display("\n2**-84 * 2**-939:");
    #10 assign a = 64'h3AB0000000000000; assign b = 64'h0540000000000000;
    #10 assign a = 64'h3ABFFFFFFFFFFFFF; assign b = 64'h054FFFFFFFFFFFFF;

    #10 $display("\n2**-83 * 2**-940:");
    #10 assign a = 64'h3AC0000000000000; assign b = 64'h0530000000000000;
    #10 assign a = 64'h3ACFFFFFFFFFFFFF; assign b = 64'h053FFFFFFFFFFFFF;

    #10 $display("\n2**-82 * 2**-941:");
    #10 assign a = 64'h3AD0000000000000; assign b = 64'h0520000000000000;
    #10 assign a = 64'h3ADFFFFFFFFFFFFF; assign b = 64'h052FFFFFFFFFFFFF;

    #10 $display("\n2**-81 * 2**-942:");
    #10 assign a = 64'h3AE0000000000000; assign b = 64'h0510000000000000;
    #10 assign a = 64'h3AEFFFFFFFFFFFFF; assign b = 64'h051FFFFFFFFFFFFF;

    #10 $display("\n2**-80 * 2**-943:");
    #10 assign a = 64'h3AF0000000000000; assign b = 64'h0500000000000000;
    #10 assign a = 64'h3AFFFFFFFFFFFFFF; assign b = 64'h050FFFFFFFFFFFFF;

    #10 $display("\n2**-79 * 2**-944:");
    #10 assign a = 64'h3B00000000000000; assign b = 64'h04F0000000000000;
    #10 assign a = 64'h3B0FFFFFFFFFFFFF; assign b = 64'h04FFFFFFFFFFFFFF;

    #10 $display("\n2**-78 * 2**-945:");
    #10 assign a = 64'h3B10000000000000; assign b = 64'h04E0000000000000;
    #10 assign a = 64'h3B1FFFFFFFFFFFFF; assign b = 64'h04EFFFFFFFFFFFFF;

    #10 $display("\n2**-77 * 2**-946:");
    #10 assign a = 64'h3B20000000000000; assign b = 64'h04D0000000000000;
    #10 assign a = 64'h3B2FFFFFFFFFFFFF; assign b = 64'h04DFFFFFFFFFFFFF;

    #10 $display("\n2**-76 * 2**-947:");
    #10 assign a = 64'h3B30000000000000; assign b = 64'h04C0000000000000;
    #10 assign a = 64'h3B3FFFFFFFFFFFFF; assign b = 64'h04CFFFFFFFFFFFFF;

    #10 $display("\n2**-75 * 2**-948:");
    #10 assign a = 64'h3B40000000000000; assign b = 64'h04B0000000000000;
    #10 assign a = 64'h3B4FFFFFFFFFFFFF; assign b = 64'h04BFFFFFFFFFFFFF;

    #10 $display("\n2**-74 * 2**-949:");
    #10 assign a = 64'h3B50000000000000; assign b = 64'h04A0000000000000;
    #10 assign a = 64'h3B5FFFFFFFFFFFFF; assign b = 64'h04AFFFFFFFFFFFFF;

    #10 $display("\n2**-73 * 2**-950:");
    #10 assign a = 64'h3B60000000000000; assign b = 64'h0490000000000000;
    #10 assign a = 64'h3B6FFFFFFFFFFFFF; assign b = 64'h049FFFFFFFFFFFFF;

    #10 $display("\n2**-72 * 2**-951:");
    #10 assign a = 64'h3B70000000000000; assign b = 64'h0480000000000000;
    #10 assign a = 64'h3B7FFFFFFFFFFFFF; assign b = 64'h048FFFFFFFFFFFFF;

    #10 $display("\n2**-71 * 2**-952:");
    #10 assign a = 64'h3B80000000000000; assign b = 64'h0470000000000000;
    #10 assign a = 64'h3B8FFFFFFFFFFFFF; assign b = 64'h047FFFFFFFFFFFFF;

    #10 $display("\n2**-70 * 2**-953:");
    #10 assign a = 64'h3B90000000000000; assign b = 64'h0460000000000000;
    #10 assign a = 64'h3B9FFFFFFFFFFFFF; assign b = 64'h046FFFFFFFFFFFFF;

    #10 $display("\n2**-69 * 2**-954:");
    #10 assign a = 64'h3BA0000000000000; assign b = 64'h0450000000000000;
    #10 assign a = 64'h3BAFFFFFFFFFFFFF; assign b = 64'h045FFFFFFFFFFFFF;

    #10 $display("\n2**-68 * 2**-955:");
    #10 assign a = 64'h3BB0000000000000; assign b = 64'h0440000000000000;
    #10 assign a = 64'h3BBFFFFFFFFFFFFF; assign b = 64'h044FFFFFFFFFFFFF;

    #10 $display("\n2**-67 * 2**-956:");
    #10 assign a = 64'h3BC0000000000000; assign b = 64'h0430000000000000;
    #10 assign a = 64'h3BCFFFFFFFFFFFFF; assign b = 64'h043FFFFFFFFFFFFF;

    #10 $display("\n2**-66 * 2**-957:");
    #10 assign a = 64'h3BD0000000000000; assign b = 64'h0420000000000000;
    #10 assign a = 64'h3BDFFFFFFFFFFFFF; assign b = 64'h042FFFFFFFFFFFFF;

    #10 $display("\n2**-65 * 2**-958:");
    #10 assign a = 64'h3BE0000000000000; assign b = 64'h0410000000000000;
    #10 assign a = 64'h3BEFFFFFFFFFFFFF; assign b = 64'h041FFFFFFFFFFFFF;

    #10 $display("\n2**-64 * 2**-959:");
    #10 assign a = 64'h3BF0000000000000; assign b = 64'h0400000000000000;
    #10 assign a = 64'h3BFFFFFFFFFFFFFF; assign b = 64'h040FFFFFFFFFFFFF;

    #10 $display("\n2**-63 * 2**-960:");
    #10 assign a = 64'h3C00000000000000; assign b = 64'h03F0000000000000;
    #10 assign a = 64'h3C0FFFFFFFFFFFFF; assign b = 64'h03FFFFFFFFFFFFFF;

    #10 $display("\n2**-62 * 2**-961:");
    #10 assign a = 64'h3C10000000000000; assign b = 64'h03E0000000000000;
    #10 assign a = 64'h3C1FFFFFFFFFFFFF; assign b = 64'h03EFFFFFFFFFFFFF;

    #10 $display("\n2**-61 * 2**-962:");
    #10 assign a = 64'h3C20000000000000; assign b = 64'h03D0000000000000;
    #10 assign a = 64'h3C2FFFFFFFFFFFFF; assign b = 64'h03DFFFFFFFFFFFFF;

    #10 $display("\n2**-60 * 2**-963:");
    #10 assign a = 64'h3C30000000000000; assign b = 64'h03C0000000000000;
    #10 assign a = 64'h3C3FFFFFFFFFFFFF; assign b = 64'h03CFFFFFFFFFFFFF;

    #10 $display("\n2**-59 * 2**-964:");
    #10 assign a = 64'h3C40000000000000; assign b = 64'h03B0000000000000;
    #10 assign a = 64'h3C4FFFFFFFFFFFFF; assign b = 64'h03BFFFFFFFFFFFFF;

    #10 $display("\n2**-58 * 2**-965:");
    #10 assign a = 64'h3C50000000000000; assign b = 64'h03A0000000000000;
    #10 assign a = 64'h3C5FFFFFFFFFFFFF; assign b = 64'h03AFFFFFFFFFFFFF;

    #10 $display("\n2**-57 * 2**-966:");
    #10 assign a = 64'h3C60000000000000; assign b = 64'h0390000000000000;
    #10 assign a = 64'h3C6FFFFFFFFFFFFF; assign b = 64'h039FFFFFFFFFFFFF;

    #10 $display("\n2**-56 * 2**-967:");
    #10 assign a = 64'h3C70000000000000; assign b = 64'h0380000000000000;
    #10 assign a = 64'h3C7FFFFFFFFFFFFF; assign b = 64'h038FFFFFFFFFFFFF;

    #10 $display("\n2**-55 * 2**-968:");
    #10 assign a = 64'h3C80000000000000; assign b = 64'h0370000000000000;
    #10 assign a = 64'h3C8FFFFFFFFFFFFF; assign b = 64'h037FFFFFFFFFFFFF;

    #10 $display("\n2**-54 * 2**-969:");
    #10 assign a = 64'h3C90000000000000; assign b = 64'h0360000000000000;
    #10 assign a = 64'h3C9FFFFFFFFFFFFF; assign b = 64'h036FFFFFFFFFFFFF;

    #10 $display("\n2**-53 * 2**-970:");
    #10 assign a = 64'h3CA0000000000000; assign b = 64'h0350000000000000;
    #10 assign a = 64'h3CAFFFFFFFFFFFFF; assign b = 64'h035FFFFFFFFFFFFF;

    #10 $display("\n2**-52 * 2**-971:");
    #10 assign a = 64'h3CB0000000000000; assign b = 64'h0340000000000000;
    #10 assign a = 64'h3CBFFFFFFFFFFFFF; assign b = 64'h034FFFFFFFFFFFFF;

    #10 $display("\n2**-51 * 2**-972:");
    #10 assign a = 64'h3CC0000000000000; assign b = 64'h0330000000000000;
    #10 assign a = 64'h3CCFFFFFFFFFFFFF; assign b = 64'h033FFFFFFFFFFFFF;

    #10 $display("\n2**-50 * 2**-973:");
    #10 assign a = 64'h3CD0000000000000; assign b = 64'h0320000000000000;
    #10 assign a = 64'h3CDFFFFFFFFFFFFF; assign b = 64'h032FFFFFFFFFFFFF;

    #10 $display("\n2**-49 * 2**-974:");
    #10 assign a = 64'h3CE0000000000000; assign b = 64'h0310000000000000;
    #10 assign a = 64'h3CEFFFFFFFFFFFFF; assign b = 64'h031FFFFFFFFFFFFF;

    #10 $display("\n2**-48 * 2**-975:");
    #10 assign a = 64'h3CF0000000000000; assign b = 64'h0300000000000000;
    #10 assign a = 64'h3CFFFFFFFFFFFFFF; assign b = 64'h030FFFFFFFFFFFFF;

    #10 $display("\n2**-47 * 2**-976:");
    #10 assign a = 64'h3D00000000000000; assign b = 64'h02F0000000000000;
    #10 assign a = 64'h3D0FFFFFFFFFFFFF; assign b = 64'h02FFFFFFFFFFFFFF;

    #10 $display("\n2**-46 * 2**-977:");
    #10 assign a = 64'h3D10000000000000; assign b = 64'h02E0000000000000;
    #10 assign a = 64'h3D1FFFFFFFFFFFFF; assign b = 64'h02EFFFFFFFFFFFFF;

    #10 $display("\n2**-45 * 2**-978:");
    #10 assign a = 64'h3D20000000000000; assign b = 64'h02D0000000000000;
    #10 assign a = 64'h3D2FFFFFFFFFFFFF; assign b = 64'h02DFFFFFFFFFFFFF;

    #10 $display("\n2**-44 * 2**-979:");
    #10 assign a = 64'h3D30000000000000; assign b = 64'h02C0000000000000;
    #10 assign a = 64'h3D3FFFFFFFFFFFFF; assign b = 64'h02CFFFFFFFFFFFFF;

    #10 $display("\n2**-43 * 2**-980:");
    #10 assign a = 64'h3D40000000000000; assign b = 64'h02B0000000000000;
    #10 assign a = 64'h3D4FFFFFFFFFFFFF; assign b = 64'h02BFFFFFFFFFFFFF;

    #10 $display("\n2**-42 * 2**-981:");
    #10 assign a = 64'h3D50000000000000; assign b = 64'h02A0000000000000;
    #10 assign a = 64'h3D5FFFFFFFFFFFFF; assign b = 64'h02AFFFFFFFFFFFFF;

    #10 $display("\n2**-41 * 2**-982:");
    #10 assign a = 64'h3D60000000000000; assign b = 64'h0290000000000000;
    #10 assign a = 64'h3D6FFFFFFFFFFFFF; assign b = 64'h029FFFFFFFFFFFFF;

    #10 $display("\n2**-40 * 2**-983:");
    #10 assign a = 64'h3D70000000000000; assign b = 64'h0280000000000000;
    #10 assign a = 64'h3D7FFFFFFFFFFFFF; assign b = 64'h028FFFFFFFFFFFFF;

    #10 $display("\n2**-39 * 2**-984:");
    #10 assign a = 64'h3D80000000000000; assign b = 64'h0270000000000000;
    #10 assign a = 64'h3D8FFFFFFFFFFFFF; assign b = 64'h027FFFFFFFFFFFFF;

    #10 $display("\n2**-38 * 2**-985:");
    #10 assign a = 64'h3D90000000000000; assign b = 64'h0260000000000000;
    #10 assign a = 64'h3D9FFFFFFFFFFFFF; assign b = 64'h026FFFFFFFFFFFFF;

    #10 $display("\n2**-37 * 2**-986:");
    #10 assign a = 64'h3DA0000000000000; assign b = 64'h0250000000000000;
    #10 assign a = 64'h3DAFFFFFFFFFFFFF; assign b = 64'h025FFFFFFFFFFFFF;

    #10 $display("\n2**-36 * 2**-987:");
    #10 assign a = 64'h3DB0000000000000; assign b = 64'h0240000000000000;
    #10 assign a = 64'h3DBFFFFFFFFFFFFF; assign b = 64'h024FFFFFFFFFFFFF;

    #10 $display("\n2**-35 * 2**-988:");
    #10 assign a = 64'h3DC0000000000000; assign b = 64'h0230000000000000;
    #10 assign a = 64'h3DCFFFFFFFFFFFFF; assign b = 64'h023FFFFFFFFFFFFF;

    #10 $display("\n2**-34 * 2**-989:");
    #10 assign a = 64'h3DD0000000000000; assign b = 64'h0220000000000000;
    #10 assign a = 64'h3DDFFFFFFFFFFFFF; assign b = 64'h022FFFFFFFFFFFFF;

    #10 $display("\n2**-33 * 2**-990:");
    #10 assign a = 64'h3DE0000000000000; assign b = 64'h0210000000000000;
    #10 assign a = 64'h3DEFFFFFFFFFFFFF; assign b = 64'h021FFFFFFFFFFFFF;

    #10 $display("\n2**-32 * 2**-991:");
    #10 assign a = 64'h3DF0000000000000; assign b = 64'h0200000000000000;
    #10 assign a = 64'h3DFFFFFFFFFFFFFF; assign b = 64'h020FFFFFFFFFFFFF;

    #10 $display("\n2**-31 * 2**-992:");
    #10 assign a = 64'h3E00000000000000; assign b = 64'h01F0000000000000;
    #10 assign a = 64'h3E0FFFFFFFFFFFFF; assign b = 64'h01FFFFFFFFFFFFFF;

    #10 $display("\n2**-30 * 2**-993:");
    #10 assign a = 64'h3E10000000000000; assign b = 64'h01E0000000000000;
    #10 assign a = 64'h3E1FFFFFFFFFFFFF; assign b = 64'h01EFFFFFFFFFFFFF;

    #10 $display("\n2**-29 * 2**-994:");
    #10 assign a = 64'h3E20000000000000; assign b = 64'h01D0000000000000;
    #10 assign a = 64'h3E2FFFFFFFFFFFFF; assign b = 64'h01DFFFFFFFFFFFFF;

    #10 $display("\n2**-28 * 2**-995:");
    #10 assign a = 64'h3E30000000000000; assign b = 64'h01C0000000000000;
    #10 assign a = 64'h3E3FFFFFFFFFFFFF; assign b = 64'h01CFFFFFFFFFFFFF;

    #10 $display("\n2**-27 * 2**-996:");
    #10 assign a = 64'h3E40000000000000; assign b = 64'h01B0000000000000;
    #10 assign a = 64'h3E4FFFFFFFFFFFFF; assign b = 64'h01BFFFFFFFFFFFFF;

    #10 $display("\n2**-26 * 2**-997:");
    #10 assign a = 64'h3E50000000000000; assign b = 64'h01A0000000000000;
    #10 assign a = 64'h3E5FFFFFFFFFFFFF; assign b = 64'h01AFFFFFFFFFFFFF;

    #10 $display("\n2**-25 * 2**-998:");
    #10 assign a = 64'h3E60000000000000; assign b = 64'h0190000000000000;
    #10 assign a = 64'h3E6FFFFFFFFFFFFF; assign b = 64'h019FFFFFFFFFFFFF;

    #10 $display("\n2**-24 * 2**-999:");
    #10 assign a = 64'h3E70000000000000; assign b = 64'h0180000000000000;
    #10 assign a = 64'h3E7FFFFFFFFFFFFF; assign b = 64'h018FFFFFFFFFFFFF;

    #10 $display("\n2**-23 * 2**-1000:");
    #10 assign a = 64'h3E80000000000000; assign b = 64'h0170000000000000;
    #10 assign a = 64'h3E8FFFFFFFFFFFFF; assign b = 64'h017FFFFFFFFFFFFF;

    #10 $display("\n2**-22 * 2**-1001:");
    #10 assign a = 64'h3E90000000000000; assign b = 64'h0160000000000000;
    #10 assign a = 64'h3E9FFFFFFFFFFFFF; assign b = 64'h016FFFFFFFFFFFFF;

    #10 $display("\n2**-21 * 2**-1002:");
    #10 assign a = 64'h3EA0000000000000; assign b = 64'h0150000000000000;
    #10 assign a = 64'h3EAFFFFFFFFFFFFF; assign b = 64'h015FFFFFFFFFFFFF;

    #10 $display("\n2**-20 * 2**-1003:");
    #10 assign a = 64'h3EB0000000000000; assign b = 64'h0140000000000000;
    #10 assign a = 64'h3EBFFFFFFFFFFFFF; assign b = 64'h014FFFFFFFFFFFFF;

    #10 $display("\n2**-19 * 2**-1004:");
    #10 assign a = 64'h3EC0000000000000; assign b = 64'h0130000000000000;
    #10 assign a = 64'h3ECFFFFFFFFFFFFF; assign b = 64'h013FFFFFFFFFFFFF;

    #10 $display("\n2**-18 * 2**-1005:");
    #10 assign a = 64'h3ED0000000000000; assign b = 64'h0120000000000000;
    #10 assign a = 64'h3EDFFFFFFFFFFFFF; assign b = 64'h012FFFFFFFFFFFFF;

    #10 $display("\n2**-17 * 2**-1006:");
    #10 assign a = 64'h3EE0000000000000; assign b = 64'h0110000000000000;
    #10 assign a = 64'h3EEFFFFFFFFFFFFF; assign b = 64'h011FFFFFFFFFFFFF;

    #10 $display("\n2**-16 * 2**-1007:");
    #10 assign a = 64'h3EF0000000000000; assign b = 64'h0100000000000000;
    #10 assign a = 64'h3EFFFFFFFFFFFFFF; assign b = 64'h010FFFFFFFFFFFFF;

    #10 $display("\n2**-15 * 2**-1008:");
    #10 assign a = 64'h3F00000000000000; assign b = 64'h00F0000000000000;
    #10 assign a = 64'h3F0FFFFFFFFFFFFF; assign b = 64'h00FFFFFFFFFFFFFF;

    #10 $display("\n2**-14 * 2**-1009:");
    #10 assign a = 64'h3F10000000000000; assign b = 64'h00E0000000000000;
    #10 assign a = 64'h3F1FFFFFFFFFFFFF; assign b = 64'h00EFFFFFFFFFFFFF;

    #10 $display("\n2**-13 * 2**-1010:");
    #10 assign a = 64'h3F20000000000000; assign b = 64'h00D0000000000000;
    #10 assign a = 64'h3F2FFFFFFFFFFFFF; assign b = 64'h00DFFFFFFFFFFFFF;

    #10 $display("\n2**-12 * 2**-1011:");
    #10 assign a = 64'h3F30000000000000; assign b = 64'h00C0000000000000;
    #10 assign a = 64'h3F3FFFFFFFFFFFFF; assign b = 64'h00CFFFFFFFFFFFFF;

    #10 $display("\n2**-11 * 2**-1012:");
    #10 assign a = 64'h3F40000000000000; assign b = 64'h00B0000000000000;
    #10 assign a = 64'h3F4FFFFFFFFFFFFF; assign b = 64'h00BFFFFFFFFFFFFF;

    #10 $display("\n2**-10 * 2**-1013:");
    #10 assign a = 64'h3F50000000000000; assign b = 64'h00A0000000000000;
    #10 assign a = 64'h3F5FFFFFFFFFFFFF; assign b = 64'h00AFFFFFFFFFFFFF;

    #10 $display("\n2**-9 * 2**-1014:");
    #10 assign a = 64'h3F60000000000000; assign b = 64'h0090000000000000;
    #10 assign a = 64'h3F6FFFFFFFFFFFFF; assign b = 64'h009FFFFFFFFFFFFF;

    #10 $display("\n2**-8 * 2**-1015:");
    #10 assign a = 64'h3F70000000000000; assign b = 64'h0080000000000000;
    #10 assign a = 64'h3F7FFFFFFFFFFFFF; assign b = 64'h008FFFFFFFFFFFFF;

    #10 $display("\n2**-7 * 2**-1016:");
    #10 assign a = 64'h3F80000000000000; assign b = 64'h0070000000000000;
    #10 assign a = 64'h3F8FFFFFFFFFFFFF; assign b = 64'h007FFFFFFFFFFFFF;

    #10 $display("\n2**-6 * 2**-1017:");
    #10 assign a = 64'h3F90000000000000; assign b = 64'h0060000000000000;
    #10 assign a = 64'h3F9FFFFFFFFFFFFF; assign b = 64'h006FFFFFFFFFFFFF;

    #10 $display("\n2**-5 * 2**-1018:");
    #10 assign a = 64'h3FA0000000000000; assign b = 64'h0050000000000000;
    #10 assign a = 64'h3FAFFFFFFFFFFFFF; assign b = 64'h005FFFFFFFFFFFFF;

    #10 $display("\n2**-4 * 2**-1019:");
    #10 assign a = 64'h3FB0000000000000; assign b = 64'h0040000000000000;
    #10 assign a = 64'h3FBFFFFFFFFFFFFF; assign b = 64'h004FFFFFFFFFFFFF;

    #10 $display("\n2**-3 * 2**-1020:");
    #10 assign a = 64'h3FC0000000000000; assign b = 64'h0030000000000000;
    #10 assign a = 64'h3FCFFFFFFFFFFFFF; assign b = 64'h003FFFFFFFFFFFFF;

    #10 $display("\n2**-2 * 2**-1021:");
    #10 assign a = 64'h3FD0000000000000; assign b = 64'h0020000000000000;
    #10 assign a = 64'h3FDFFFFFFFFFFFFF; assign b = 64'h002FFFFFFFFFFFFF;

    #10 $display("\n2**-1 * 2**-1022:");
    #10 assign a = 64'h3FE0000000000000; assign b = 64'h0010000000000000;
    #10 assign a = 64'h3FEFFFFFFFFFFFFF; assign b = 64'h001FFFFFFFFFFFFF;

    #10 $display("\n2**0 * 2**-1023:");
    #10 assign a = 64'h3FF0000000000000; assign b = 64'h0008000000000000;
    #10 assign a = 64'h3FFFFFFFFFFFFFFF; assign b = 64'h000FFFFFFFFFFFFF;

    #10 $display("\n2**1 * 2**-1024:");
    #10 assign a = 64'h4000000000000000; assign b = 64'h0004000000000000;
    #10 assign a = 64'h400FFFFFFFFFFFFF; assign b = 64'h0007FFFFFFFFFFFF;

    #10 $display("\n2**2 * 2**-1025:");
    #10 assign a = 64'h4010000000000000; assign b = 64'h0002000000000000;
    #10 assign a = 64'h401FFFFFFFFFFFFF; assign b = 64'h0003FFFFFFFFFFFF;

    #10 $display("\n2**3 * 2**-1026:");
    #10 assign a = 64'h4020000000000000; assign b = 64'h0001000000000000;
    #10 assign a = 64'h402FFFFFFFFFFFFF; assign b = 64'h0001FFFFFFFFFFFF;

    #10 $display("\n2**4 * 2**-1027:");
    #10 assign a = 64'h4030000000000000; assign b = 64'h0000800000000000;
    #10 assign a = 64'h403FFFFFFFFFFFFF; assign b = 64'h0000FFFFFFFFFFFF;

    #10 $display("\n2**5 * 2**-1028:");
    #10 assign a = 64'h4040000000000000; assign b = 64'h0000400000000000;
    #10 assign a = 64'h404FFFFFFFFFFFFF; assign b = 64'h00007FFFFFFFFFFF;

    #10 $display("\n2**6 * 2**-1029:");
    #10 assign a = 64'h4050000000000000; assign b = 64'h0000200000000000;
    #10 assign a = 64'h405FFFFFFFFFFFFF; assign b = 64'h00003FFFFFFFFFFF;

    #10 $display("\n2**7 * 2**-1030:");
    #10 assign a = 64'h4060000000000000; assign b = 64'h0000100000000000;
    #10 assign a = 64'h406FFFFFFFFFFFFF; assign b = 64'h00001FFFFFFFFFFF;

    #10 $display("\n2**8 * 2**-1031:");
    #10 assign a = 64'h4070000000000000; assign b = 64'h0000080000000000;
    #10 assign a = 64'h407FFFFFFFFFFFFF; assign b = 64'h00000FFFFFFFFFFF;

    #10 $display("\n2**9 * 2**-1032:");
    #10 assign a = 64'h4080000000000000; assign b = 64'h0000040000000000;
    #10 assign a = 64'h408FFFFFFFFFFFFF; assign b = 64'h000007FFFFFFFFFF;

    #10 $display("\n2**10 * 2**-1033:");
    #10 assign a = 64'h4090000000000000; assign b = 64'h0000020000000000;
    #10 assign a = 64'h409FFFFFFFFFFFFF; assign b = 64'h000003FFFFFFFFFF;

    #10 $display("\n2**11 * 2**-1034:");
    #10 assign a = 64'h40A0000000000000; assign b = 64'h0000010000000000;
    #10 assign a = 64'h40AFFFFFFFFFFFFF; assign b = 64'h000001FFFFFFFFFF;

    #10 $display("\n2**12 * 2**-1035:");
    #10 assign a = 64'h40B0000000000000; assign b = 64'h0000008000000000;
    #10 assign a = 64'h40BFFFFFFFFFFFFF; assign b = 64'h000000FFFFFFFFFF;

    #10 $display("\n2**13 * 2**-1036:");
    #10 assign a = 64'h40C0000000000000; assign b = 64'h0000004000000000;
    #10 assign a = 64'h40CFFFFFFFFFFFFF; assign b = 64'h0000007FFFFFFFFF;

    #10 $display("\n2**14 * 2**-1037:");
    #10 assign a = 64'h40D0000000000000; assign b = 64'h0000002000000000;
    #10 assign a = 64'h40DFFFFFFFFFFFFF; assign b = 64'h0000003FFFFFFFFF;

    #10 $display("\n2**15 * 2**-1038:");
    #10 assign a = 64'h40E0000000000000; assign b = 64'h0000001000000000;
    #10 assign a = 64'h40EFFFFFFFFFFFFF; assign b = 64'h0000001FFFFFFFFF;

    #10 $display("\n2**16 * 2**-1039:");
    #10 assign a = 64'h40F0000000000000; assign b = 64'h0000000800000000;
    #10 assign a = 64'h40FFFFFFFFFFFFFF; assign b = 64'h0000000FFFFFFFFF;

    #10 $display("\n2**17 * 2**-1040:");
    #10 assign a = 64'h4100000000000000; assign b = 64'h0000000400000000;
    #10 assign a = 64'h410FFFFFFFFFFFFF; assign b = 64'h00000007FFFFFFFF;

    #10 $display("\n2**18 * 2**-1041:");
    #10 assign a = 64'h4110000000000000; assign b = 64'h0000000200000000;
    #10 assign a = 64'h411FFFFFFFFFFFFF; assign b = 64'h00000003FFFFFFFF;

    #10 $display("\n2**19 * 2**-1042:");
    #10 assign a = 64'h4120000000000000; assign b = 64'h0000000100000000;
    #10 assign a = 64'h412FFFFFFFFFFFFF; assign b = 64'h00000001FFFFFFFF;

    #10 $display("\n2**20 * 2**-1043:");
    #10 assign a = 64'h4130000000000000; assign b = 64'h0000000080000000;
    #10 assign a = 64'h413FFFFFFFFFFFFF; assign b = 64'h00000000FFFFFFFF;

    #10 $display("\n2**21 * 2**-1044:");
    #10 assign a = 64'h4140000000000000; assign b = 64'h0000000040000000;
    #10 assign a = 64'h414FFFFFFFFFFFFF; assign b = 64'h000000007FFFFFFF;

    #10 $display("\n2**22 * 2**-1045:");
    #10 assign a = 64'h4150000000000000; assign b = 64'h0000000020000000;
    #10 assign a = 64'h415FFFFFFFFFFFFF; assign b = 64'h000000003FFFFFFF;

    #10 $display("\n2**23 * 2**-1046:");
    #10 assign a = 64'h4160000000000000; assign b = 64'h0000000010000000;
    #10 assign a = 64'h416FFFFFFFFFFFFF; assign b = 64'h000000001FFFFFFF;

    #10 $display("\n2**24 * 2**-1047:");
    #10 assign a = 64'h4170000000000000; assign b = 64'h0000000008000000;
    #10 assign a = 64'h417FFFFFFFFFFFFF; assign b = 64'h000000000FFFFFFF;

    #10 $display("\n2**25 * 2**-1048:");
    #10 assign a = 64'h4180000000000000; assign b = 64'h0000000004000000;
    #10 assign a = 64'h418FFFFFFFFFFFFF; assign b = 64'h0000000007FFFFFF;

    #10 $display("\n2**26 * 2**-1049:");
    #10 assign a = 64'h4190000000000000; assign b = 64'h0000000002000000;
    #10 assign a = 64'h419FFFFFFFFFFFFF; assign b = 64'h0000000003FFFFFF;

    #10 $display("\n2**27 * 2**-1050:");
    #10 assign a = 64'h41A0000000000000; assign b = 64'h0000000001000000;
    #10 assign a = 64'h41AFFFFFFFFFFFFF; assign b = 64'h0000000001FFFFFF;

    #10 $display("\n2**28 * 2**-1051:");
    #10 assign a = 64'h41B0000000000000; assign b = 64'h0000000000800000;
    #10 assign a = 64'h41BFFFFFFFFFFFFF; assign b = 64'h0000000000FFFFFF;

    #10 $display("\n2**29 * 2**-1052:");
    #10 assign a = 64'h41C0000000000000; assign b = 64'h0000000000400000;
    #10 assign a = 64'h41CFFFFFFFFFFFFF; assign b = 64'h00000000007FFFFF;

    #10 $display("\n2**30 * 2**-1053:");
    #10 assign a = 64'h41D0000000000000; assign b = 64'h0000000000200000;
    #10 assign a = 64'h41DFFFFFFFFFFFFF; assign b = 64'h00000000003FFFFF;

    #10 $display("\n2**31 * 2**-1054:");
    #10 assign a = 64'h41E0000000000000; assign b = 64'h0000000000100000;
    #10 assign a = 64'h41EFFFFFFFFFFFFF; assign b = 64'h00000000001FFFFF;

    #10 $display("\n2**32 * 2**-1055:");
    #10 assign a = 64'h41F0000000000000; assign b = 64'h0000000000080000;
    #10 assign a = 64'h41FFFFFFFFFFFFFF; assign b = 64'h00000000000FFFFF;

    #10 $display("\n2**33 * 2**-1056:");
    #10 assign a = 64'h4200000000000000; assign b = 64'h0000000000040000;
    #10 assign a = 64'h420FFFFFFFFFFFFF; assign b = 64'h000000000007FFFF;

    #10 $display("\n2**34 * 2**-1057:");
    #10 assign a = 64'h4210000000000000; assign b = 64'h0000000000020000;
    #10 assign a = 64'h421FFFFFFFFFFFFF; assign b = 64'h000000000003FFFF;

    #10 $display("\n2**35 * 2**-1058:");
    #10 assign a = 64'h4220000000000000; assign b = 64'h0000000000010000;
    #10 assign a = 64'h422FFFFFFFFFFFFF; assign b = 64'h000000000001FFFF;

    #10 $display("\n2**36 * 2**-1059:");
    #10 assign a = 64'h4230000000000000; assign b = 64'h0000000000008000;
    #10 assign a = 64'h423FFFFFFFFFFFFF; assign b = 64'h000000000000FFFF;

    #10 $display("\n2**37 * 2**-1060:");
    #10 assign a = 64'h4240000000000000; assign b = 64'h0000000000004000;
    #10 assign a = 64'h424FFFFFFFFFFFFF; assign b = 64'h0000000000007FFF;

    #10 $display("\n2**38 * 2**-1061:");
    #10 assign a = 64'h4250000000000000; assign b = 64'h0000000000002000;
    #10 assign a = 64'h425FFFFFFFFFFFFF; assign b = 64'h0000000000003FFF;

    #10 $display("\n2**39 * 2**-1062:");
    #10 assign a = 64'h4260000000000000; assign b = 64'h0000000000001000;
    #10 assign a = 64'h426FFFFFFFFFFFFF; assign b = 64'h0000000000001FFF;

    #10 $display("\n2**40 * 2**-1063:");
    #10 assign a = 64'h4270000000000000; assign b = 64'h0000000000000800;
    #10 assign a = 64'h427FFFFFFFFFFFFF; assign b = 64'h0000000000000FFF;

    #10 $display("\n2**41 * 2**-1064:");
    #10 assign a = 64'h4280000000000000; assign b = 64'h0000000000000400;
    #10 assign a = 64'h428FFFFFFFFFFFFF; assign b = 64'h00000000000007FF;

    #10 $display("\n2**42 * 2**-1065:");
    #10 assign a = 64'h4290000000000000; assign b = 64'h0000000000000200;
    #10 assign a = 64'h429FFFFFFFFFFFFF; assign b = 64'h00000000000003FF;

    #10 $display("\n2**43 * 2**-1066:");
    #10 assign a = 64'h42A0000000000000; assign b = 64'h0000000000000100;
    #10 assign a = 64'h42AFFFFFFFFFFFFF; assign b = 64'h00000000000001FF;

    #10 $display("\n2**44 * 2**-1067:");
    #10 assign a = 64'h42B0000000000000; assign b = 64'h0000000000000080;
    #10 assign a = 64'h42BFFFFFFFFFFFFF; assign b = 64'h00000000000000FF;

    #10 $display("\n2**45 * 2**-1068:");
    #10 assign a = 64'h42C0000000000000; assign b = 64'h0000000000000040;
    #10 assign a = 64'h42CFFFFFFFFFFFFF; assign b = 64'h000000000000007F;

    #10 $display("\n2**46 * 2**-1069:");
    #10 assign a = 64'h42D0000000000000; assign b = 64'h0000000000000020;
    #10 assign a = 64'h42DFFFFFFFFFFFFF; assign b = 64'h000000000000003F;

    #10 $display("\n2**47 * 2**-1070:");
    #10 assign a = 64'h42E0000000000000; assign b = 64'h0000000000000010;
    #10 assign a = 64'h42EFFFFFFFFFFFFF; assign b = 64'h000000000000001F;

    #10 $display("\n2**48 * 2**-1071:");
    #10 assign a = 64'h42F0000000000000; assign b = 64'h0000000000000008;
    #10 assign a = 64'h42FFFFFFFFFFFFFF; assign b = 64'h000000000000000F;

    #10 $display("\n2**49 * 2**-1072:");
    #10 assign a = 64'h4300000000000000; assign b = 64'h0000000000000004;
    #10 assign a = 64'h430FFFFFFFFFFFFF; assign b = 64'h0000000000000007;

    #10 $display("\n2**50 * 2**-1073:");
    #10 assign a = 64'h4310000000000000; assign b = 64'h0000000000000002;
    #10 assign a = 64'h431FFFFFFFFFFFFF; assign b = 64'h0000000000000003;

    #10 $display("\n2**51 * 2**-1074:");
    #10 assign a = 64'h4320000000000000; assign b = 64'h0000000000000001;
    #10 assign a = 64'h432FFFFFFFFFFFFF; assign b = 64'h0000000000000001;

    #10 $display("\n2**-1074 * 2**-1:");
    #10 assign a = 64'h0000000000000001; assign b = 64'h3FE0000000000000;
    #10 assign a = 64'h0000000000000001; assign b = 64'h3FEFFFFFFFFFFFFF;

    #10 $display("\n2**-1073 * 2**-2:");
    #10 assign a = 64'h0000000000000002; assign b = 64'h3FD0000000000000;
    #10 assign a = 64'h0000000000000003; assign b = 64'h3FDFFFFFFFFFFFFF;

    #10 $display("\n2**-1072 * 2**-3:");
    #10 assign a = 64'h0000000000000004; assign b = 64'h3FC0000000000000;
    #10 assign a = 64'h0000000000000007; assign b = 64'h3FCFFFFFFFFFFFFF;

    #10 $display("\n2**-1071 * 2**-4:");
    #10 assign a = 64'h0000000000000008; assign b = 64'h3FB0000000000000;
    #10 assign a = 64'h000000000000000F; assign b = 64'h3FBFFFFFFFFFFFFF;

    #10 $display("\n2**-1070 * 2**-5:");
    #10 assign a = 64'h0000000000000010; assign b = 64'h3FA0000000000000;
    #10 assign a = 64'h000000000000001F; assign b = 64'h3FAFFFFFFFFFFFFF;

    #10 $display("\n2**-1069 * 2**-6:");
    #10 assign a = 64'h0000000000000020; assign b = 64'h3F90000000000000;
    #10 assign a = 64'h000000000000003F; assign b = 64'h3F9FFFFFFFFFFFFF;

    #10 $display("\n2**-1068 * 2**-7:");
    #10 assign a = 64'h0000000000000040; assign b = 64'h3F80000000000000;
    #10 assign a = 64'h000000000000007F; assign b = 64'h3F8FFFFFFFFFFFFF;

    #10 $display("\n2**-1067 * 2**-8:");
    #10 assign a = 64'h0000000000000080; assign b = 64'h3F70000000000000;
    #10 assign a = 64'h00000000000000FF; assign b = 64'h3F7FFFFFFFFFFFFF;

    #10 $display("\n2**-1066 * 2**-9:");
    #10 assign a = 64'h0000000000000100; assign b = 64'h3F60000000000000;
    #10 assign a = 64'h00000000000001FF; assign b = 64'h3F6FFFFFFFFFFFFF;

    #10 $display("\n2**-1065 * 2**-10:");
    #10 assign a = 64'h0000000000000200; assign b = 64'h3F50000000000000;
    #10 assign a = 64'h00000000000003FF; assign b = 64'h3F5FFFFFFFFFFFFF;

    #10 $display("\n2**-1064 * 2**-11:");
    #10 assign a = 64'h0000000000000400; assign b = 64'h3F40000000000000;
    #10 assign a = 64'h00000000000007FF; assign b = 64'h3F4FFFFFFFFFFFFF;

    #10 $display("\n2**-1063 * 2**-12:");
    #10 assign a = 64'h0000000000000800; assign b = 64'h3F30000000000000;
    #10 assign a = 64'h0000000000000FFF; assign b = 64'h3F3FFFFFFFFFFFFF;

    #10 $display("\n2**-1062 * 2**-13:");
    #10 assign a = 64'h0000000000001000; assign b = 64'h3F20000000000000;
    #10 assign a = 64'h0000000000001FFF; assign b = 64'h3F2FFFFFFFFFFFFF;

    #10 $display("\n2**-1061 * 2**-14:");
    #10 assign a = 64'h0000000000002000; assign b = 64'h3F10000000000000;
    #10 assign a = 64'h0000000000003FFF; assign b = 64'h3F1FFFFFFFFFFFFF;

    #10 $display("\n2**-1060 * 2**-15:");
    #10 assign a = 64'h0000000000004000; assign b = 64'h3F00000000000000;
    #10 assign a = 64'h0000000000007FFF; assign b = 64'h3F0FFFFFFFFFFFFF;

    #10 $display("\n2**-1059 * 2**-16:");
    #10 assign a = 64'h0000000000008000; assign b = 64'h3EF0000000000000;
    #10 assign a = 64'h000000000000FFFF; assign b = 64'h3EFFFFFFFFFFFFFF;

    #10 $display("\n2**-1058 * 2**-17:");
    #10 assign a = 64'h0000000000010000; assign b = 64'h3EE0000000000000;
    #10 assign a = 64'h000000000001FFFF; assign b = 64'h3EEFFFFFFFFFFFFF;

    #10 $display("\n2**-1057 * 2**-18:");
    #10 assign a = 64'h0000000000020000; assign b = 64'h3ED0000000000000;
    #10 assign a = 64'h000000000003FFFF; assign b = 64'h3EDFFFFFFFFFFFFF;

    #10 $display("\n2**-1056 * 2**-19:");
    #10 assign a = 64'h0000000000040000; assign b = 64'h3EC0000000000000;
    #10 assign a = 64'h000000000007FFFF; assign b = 64'h3ECFFFFFFFFFFFFF;

    #10 $display("\n2**-1055 * 2**-20:");
    #10 assign a = 64'h0000000000080000; assign b = 64'h3EB0000000000000;
    #10 assign a = 64'h00000000000FFFFF; assign b = 64'h3EBFFFFFFFFFFFFF;

    #10 $display("\n2**-1054 * 2**-21:");
    #10 assign a = 64'h0000000000100000; assign b = 64'h3EA0000000000000;
    #10 assign a = 64'h00000000001FFFFF; assign b = 64'h3EAFFFFFFFFFFFFF;

    #10 $display("\n2**-1053 * 2**-22:");
    #10 assign a = 64'h0000000000200000; assign b = 64'h3E90000000000000;
    #10 assign a = 64'h00000000003FFFFF; assign b = 64'h3E9FFFFFFFFFFFFF;

    #10 $display("\n2**-1052 * 2**-23:");
    #10 assign a = 64'h0000000000400000; assign b = 64'h3E80000000000000;
    #10 assign a = 64'h00000000007FFFFF; assign b = 64'h3E8FFFFFFFFFFFFF;

    #10 $display("\n2**-1051 * 2**-24:");
    #10 assign a = 64'h0000000000800000; assign b = 64'h3E70000000000000;
    #10 assign a = 64'h0000000000FFFFFF; assign b = 64'h3E7FFFFFFFFFFFFF;

    #10 $display("\n2**-1050 * 2**-25:");
    #10 assign a = 64'h0000000001000000; assign b = 64'h3E60000000000000;
    #10 assign a = 64'h0000000001FFFFFF; assign b = 64'h3E6FFFFFFFFFFFFF;

    #10 $display("\n2**-1049 * 2**-26:");
    #10 assign a = 64'h0000000002000000; assign b = 64'h3E50000000000000;
    #10 assign a = 64'h0000000003FFFFFF; assign b = 64'h3E5FFFFFFFFFFFFF;

    #10 $display("\n2**-1048 * 2**-27:");
    #10 assign a = 64'h0000000004000000; assign b = 64'h3E40000000000000;
    #10 assign a = 64'h0000000007FFFFFF; assign b = 64'h3E4FFFFFFFFFFFFF;

    #10 $display("\n2**-1047 * 2**-28:");
    #10 assign a = 64'h0000000008000000; assign b = 64'h3E30000000000000;
    #10 assign a = 64'h000000000FFFFFFF; assign b = 64'h3E3FFFFFFFFFFFFF;

    #10 $display("\n2**-1046 * 2**-29:");
    #10 assign a = 64'h0000000010000000; assign b = 64'h3E20000000000000;
    #10 assign a = 64'h000000001FFFFFFF; assign b = 64'h3E2FFFFFFFFFFFFF;

    #10 $display("\n2**-1045 * 2**-30:");
    #10 assign a = 64'h0000000020000000; assign b = 64'h3E10000000000000;
    #10 assign a = 64'h000000003FFFFFFF; assign b = 64'h3E1FFFFFFFFFFFFF;

    #10 $display("\n2**-1044 * 2**-31:");
    #10 assign a = 64'h0000000040000000; assign b = 64'h3E00000000000000;
    #10 assign a = 64'h000000007FFFFFFF; assign b = 64'h3E0FFFFFFFFFFFFF;

    #10 $display("\n2**-1043 * 2**-32:");
    #10 assign a = 64'h0000000080000000; assign b = 64'h3DF0000000000000;
    #10 assign a = 64'h00000000FFFFFFFF; assign b = 64'h3DFFFFFFFFFFFFFF;

    #10 $display("\n2**-1042 * 2**-33:");
    #10 assign a = 64'h0000000100000000; assign b = 64'h3DE0000000000000;
    #10 assign a = 64'h00000001FFFFFFFF; assign b = 64'h3DEFFFFFFFFFFFFF;

    #10 $display("\n2**-1041 * 2**-34:");
    #10 assign a = 64'h0000000200000000; assign b = 64'h3DD0000000000000;
    #10 assign a = 64'h00000003FFFFFFFF; assign b = 64'h3DDFFFFFFFFFFFFF;

    #10 $display("\n2**-1040 * 2**-35:");
    #10 assign a = 64'h0000000400000000; assign b = 64'h3DC0000000000000;
    #10 assign a = 64'h00000007FFFFFFFF; assign b = 64'h3DCFFFFFFFFFFFFF;

    #10 $display("\n2**-1039 * 2**-36:");
    #10 assign a = 64'h0000000800000000; assign b = 64'h3DB0000000000000;
    #10 assign a = 64'h0000000FFFFFFFFF; assign b = 64'h3DBFFFFFFFFFFFFF;

    #10 $display("\n2**-1038 * 2**-37:");
    #10 assign a = 64'h0000001000000000; assign b = 64'h3DA0000000000000;
    #10 assign a = 64'h0000001FFFFFFFFF; assign b = 64'h3DAFFFFFFFFFFFFF;

    #10 $display("\n2**-1037 * 2**-38:");
    #10 assign a = 64'h0000002000000000; assign b = 64'h3D90000000000000;
    #10 assign a = 64'h0000003FFFFFFFFF; assign b = 64'h3D9FFFFFFFFFFFFF;

    #10 $display("\n2**-1036 * 2**-39:");
    #10 assign a = 64'h0000004000000000; assign b = 64'h3D80000000000000;
    #10 assign a = 64'h0000007FFFFFFFFF; assign b = 64'h3D8FFFFFFFFFFFFF;

    #10 $display("\n2**-1035 * 2**-40:");
    #10 assign a = 64'h0000008000000000; assign b = 64'h3D70000000000000;
    #10 assign a = 64'h000000FFFFFFFFFF; assign b = 64'h3D7FFFFFFFFFFFFF;

    #10 $display("\n2**-1034 * 2**-41:");
    #10 assign a = 64'h0000010000000000; assign b = 64'h3D60000000000000;
    #10 assign a = 64'h000001FFFFFFFFFF; assign b = 64'h3D6FFFFFFFFFFFFF;

    #10 $display("\n2**-1033 * 2**-42:");
    #10 assign a = 64'h0000020000000000; assign b = 64'h3D50000000000000;
    #10 assign a = 64'h000003FFFFFFFFFF; assign b = 64'h3D5FFFFFFFFFFFFF;

    #10 $display("\n2**-1032 * 2**-43:");
    #10 assign a = 64'h0000040000000000; assign b = 64'h3D40000000000000;
    #10 assign a = 64'h000007FFFFFFFFFF; assign b = 64'h3D4FFFFFFFFFFFFF;

    #10 $display("\n2**-1031 * 2**-44:");
    #10 assign a = 64'h0000080000000000; assign b = 64'h3D30000000000000;
    #10 assign a = 64'h00000FFFFFFFFFFF; assign b = 64'h3D3FFFFFFFFFFFFF;

    #10 $display("\n2**-1030 * 2**-45:");
    #10 assign a = 64'h0000100000000000; assign b = 64'h3D20000000000000;
    #10 assign a = 64'h00001FFFFFFFFFFF; assign b = 64'h3D2FFFFFFFFFFFFF;

    #10 $display("\n2**-1029 * 2**-46:");
    #10 assign a = 64'h0000200000000000; assign b = 64'h3D10000000000000;
    #10 assign a = 64'h00003FFFFFFFFFFF; assign b = 64'h3D1FFFFFFFFFFFFF;

    #10 $display("\n2**-1028 * 2**-47:");
    #10 assign a = 64'h0000400000000000; assign b = 64'h3D00000000000000;
    #10 assign a = 64'h00007FFFFFFFFFFF; assign b = 64'h3D0FFFFFFFFFFFFF;

    #10 $display("\n2**-1027 * 2**-48:");
    #10 assign a = 64'h0000800000000000; assign b = 64'h3CF0000000000000;
    #10 assign a = 64'h0000FFFFFFFFFFFF; assign b = 64'h3CFFFFFFFFFFFFFF;

    #10 $display("\n2**-1026 * 2**-49:");
    #10 assign a = 64'h0001000000000000; assign b = 64'h3CE0000000000000;
    #10 assign a = 64'h0001FFFFFFFFFFFF; assign b = 64'h3CEFFFFFFFFFFFFF;

    #10 $display("\n2**-1025 * 2**-50:");
    #10 assign a = 64'h0002000000000000; assign b = 64'h3CD0000000000000;
    #10 assign a = 64'h0003FFFFFFFFFFFF; assign b = 64'h3CDFFFFFFFFFFFFF;

    #10 $display("\n2**-1024 * 2**-51:");
    #10 assign a = 64'h0004000000000000; assign b = 64'h3CC0000000000000;
    #10 assign a = 64'h0007FFFFFFFFFFFF; assign b = 64'h3CCFFFFFFFFFFFFF;

    #10 $display("\n2**-1023 * 2**-52:");
    #10 assign a = 64'h0008000000000000; assign b = 64'h3CB0000000000000;
    #10 assign a = 64'h000FFFFFFFFFFFFF; assign b = 64'h3CBFFFFFFFFFFFFF;

    #10 $display("\n2**-1022 * 2**-53:");
    #10 assign a = 64'h0010000000000000; assign b = 64'h3CA0000000000000;
    #10 assign a = 64'h001FFFFFFFFFFFFF; assign b = 64'h3CAFFFFFFFFFFFFF;

    #10 $display("\n2**-1021 * 2**-54:");
    #10 assign a = 64'h0020000000000000; assign b = 64'h3C90000000000000;
    #10 assign a = 64'h002FFFFFFFFFFFFF; assign b = 64'h3C9FFFFFFFFFFFFF;

    #10 $display("\n2**-1020 * 2**-55:");
    #10 assign a = 64'h0030000000000000; assign b = 64'h3C80000000000000;
    #10 assign a = 64'h003FFFFFFFFFFFFF; assign b = 64'h3C8FFFFFFFFFFFFF;

    #10 $display("\n2**-1019 * 2**-56:");
    #10 assign a = 64'h0040000000000000; assign b = 64'h3C70000000000000;
    #10 assign a = 64'h004FFFFFFFFFFFFF; assign b = 64'h3C7FFFFFFFFFFFFF;

    #10 $display("\n2**-1018 * 2**-57:");
    #10 assign a = 64'h0050000000000000; assign b = 64'h3C60000000000000;
    #10 assign a = 64'h005FFFFFFFFFFFFF; assign b = 64'h3C6FFFFFFFFFFFFF;

    #10 $display("\n2**-1017 * 2**-58:");
    #10 assign a = 64'h0060000000000000; assign b = 64'h3C50000000000000;
    #10 assign a = 64'h006FFFFFFFFFFFFF; assign b = 64'h3C5FFFFFFFFFFFFF;

    #10 $display("\n2**-1016 * 2**-59:");
    #10 assign a = 64'h0070000000000000; assign b = 64'h3C40000000000000;
    #10 assign a = 64'h007FFFFFFFFFFFFF; assign b = 64'h3C4FFFFFFFFFFFFF;

    #10 $display("\n2**-1015 * 2**-60:");
    #10 assign a = 64'h0080000000000000; assign b = 64'h3C30000000000000;
    #10 assign a = 64'h008FFFFFFFFFFFFF; assign b = 64'h3C3FFFFFFFFFFFFF;

    #10 $display("\n2**-1014 * 2**-61:");
    #10 assign a = 64'h0090000000000000; assign b = 64'h3C20000000000000;
    #10 assign a = 64'h009FFFFFFFFFFFFF; assign b = 64'h3C2FFFFFFFFFFFFF;

    #10 $display("\n2**-1013 * 2**-62:");
    #10 assign a = 64'h00A0000000000000; assign b = 64'h3C10000000000000;
    #10 assign a = 64'h00AFFFFFFFFFFFFF; assign b = 64'h3C1FFFFFFFFFFFFF;

    #10 $display("\n2**-1012 * 2**-63:");
    #10 assign a = 64'h00B0000000000000; assign b = 64'h3C00000000000000;
    #10 assign a = 64'h00BFFFFFFFFFFFFF; assign b = 64'h3C0FFFFFFFFFFFFF;

    #10 $display("\n2**-1011 * 2**-64:");
    #10 assign a = 64'h00C0000000000000; assign b = 64'h3BF0000000000000;
    #10 assign a = 64'h00CFFFFFFFFFFFFF; assign b = 64'h3BFFFFFFFFFFFFFF;

    #10 $display("\n2**-1010 * 2**-65:");
    #10 assign a = 64'h00D0000000000000; assign b = 64'h3BE0000000000000;
    #10 assign a = 64'h00DFFFFFFFFFFFFF; assign b = 64'h3BEFFFFFFFFFFFFF;

    #10 $display("\n2**-1009 * 2**-66:");
    #10 assign a = 64'h00E0000000000000; assign b = 64'h3BD0000000000000;
    #10 assign a = 64'h00EFFFFFFFFFFFFF; assign b = 64'h3BDFFFFFFFFFFFFF;

    #10 $display("\n2**-1008 * 2**-67:");
    #10 assign a = 64'h00F0000000000000; assign b = 64'h3BC0000000000000;
    #10 assign a = 64'h00FFFFFFFFFFFFFF; assign b = 64'h3BCFFFFFFFFFFFFF;

    #10 $display("\n2**-1007 * 2**-68:");
    #10 assign a = 64'h0100000000000000; assign b = 64'h3BB0000000000000;
    #10 assign a = 64'h010FFFFFFFFFFFFF; assign b = 64'h3BBFFFFFFFFFFFFF;

    #10 $display("\n2**-1006 * 2**-69:");
    #10 assign a = 64'h0110000000000000; assign b = 64'h3BA0000000000000;
    #10 assign a = 64'h011FFFFFFFFFFFFF; assign b = 64'h3BAFFFFFFFFFFFFF;

    #10 $display("\n2**-1005 * 2**-70:");
    #10 assign a = 64'h0120000000000000; assign b = 64'h3B90000000000000;
    #10 assign a = 64'h012FFFFFFFFFFFFF; assign b = 64'h3B9FFFFFFFFFFFFF;

    #10 $display("\n2**-1004 * 2**-71:");
    #10 assign a = 64'h0130000000000000; assign b = 64'h3B80000000000000;
    #10 assign a = 64'h013FFFFFFFFFFFFF; assign b = 64'h3B8FFFFFFFFFFFFF;

    #10 $display("\n2**-1003 * 2**-72:");
    #10 assign a = 64'h0140000000000000; assign b = 64'h3B70000000000000;
    #10 assign a = 64'h014FFFFFFFFFFFFF; assign b = 64'h3B7FFFFFFFFFFFFF;

    #10 $display("\n2**-1002 * 2**-73:");
    #10 assign a = 64'h0150000000000000; assign b = 64'h3B60000000000000;
    #10 assign a = 64'h015FFFFFFFFFFFFF; assign b = 64'h3B6FFFFFFFFFFFFF;

    #10 $display("\n2**-1001 * 2**-74:");
    #10 assign a = 64'h0160000000000000; assign b = 64'h3B50000000000000;
    #10 assign a = 64'h016FFFFFFFFFFFFF; assign b = 64'h3B5FFFFFFFFFFFFF;

    #10 $display("\n2**-1000 * 2**-75:");
    #10 assign a = 64'h0170000000000000; assign b = 64'h3B40000000000000;
    #10 assign a = 64'h017FFFFFFFFFFFFF; assign b = 64'h3B4FFFFFFFFFFFFF;

    #10 $display("\n2**-999 * 2**-76:");
    #10 assign a = 64'h0180000000000000; assign b = 64'h3B30000000000000;
    #10 assign a = 64'h018FFFFFFFFFFFFF; assign b = 64'h3B3FFFFFFFFFFFFF;

    #10 $display("\n2**-998 * 2**-77:");
    #10 assign a = 64'h0190000000000000; assign b = 64'h3B20000000000000;
    #10 assign a = 64'h019FFFFFFFFFFFFF; assign b = 64'h3B2FFFFFFFFFFFFF;

    #10 $display("\n2**-997 * 2**-78:");
    #10 assign a = 64'h01A0000000000000; assign b = 64'h3B10000000000000;
    #10 assign a = 64'h01AFFFFFFFFFFFFF; assign b = 64'h3B1FFFFFFFFFFFFF;

    #10 $display("\n2**-996 * 2**-79:");
    #10 assign a = 64'h01B0000000000000; assign b = 64'h3B00000000000000;
    #10 assign a = 64'h01BFFFFFFFFFFFFF; assign b = 64'h3B0FFFFFFFFFFFFF;

    #10 $display("\n2**-995 * 2**-80:");
    #10 assign a = 64'h01C0000000000000; assign b = 64'h3AF0000000000000;
    #10 assign a = 64'h01CFFFFFFFFFFFFF; assign b = 64'h3AFFFFFFFFFFFFFF;

    #10 $display("\n2**-994 * 2**-81:");
    #10 assign a = 64'h01D0000000000000; assign b = 64'h3AE0000000000000;
    #10 assign a = 64'h01DFFFFFFFFFFFFF; assign b = 64'h3AEFFFFFFFFFFFFF;

    #10 $display("\n2**-993 * 2**-82:");
    #10 assign a = 64'h01E0000000000000; assign b = 64'h3AD0000000000000;
    #10 assign a = 64'h01EFFFFFFFFFFFFF; assign b = 64'h3ADFFFFFFFFFFFFF;

    #10 $display("\n2**-992 * 2**-83:");
    #10 assign a = 64'h01F0000000000000; assign b = 64'h3AC0000000000000;
    #10 assign a = 64'h01FFFFFFFFFFFFFF; assign b = 64'h3ACFFFFFFFFFFFFF;

    #10 $display("\n2**-991 * 2**-84:");
    #10 assign a = 64'h0200000000000000; assign b = 64'h3AB0000000000000;
    #10 assign a = 64'h020FFFFFFFFFFFFF; assign b = 64'h3ABFFFFFFFFFFFFF;

    #10 $display("\n2**-990 * 2**-85:");
    #10 assign a = 64'h0210000000000000; assign b = 64'h3AA0000000000000;
    #10 assign a = 64'h021FFFFFFFFFFFFF; assign b = 64'h3AAFFFFFFFFFFFFF;

    #10 $display("\n2**-989 * 2**-86:");
    #10 assign a = 64'h0220000000000000; assign b = 64'h3A90000000000000;
    #10 assign a = 64'h022FFFFFFFFFFFFF; assign b = 64'h3A9FFFFFFFFFFFFF;

    #10 $display("\n2**-988 * 2**-87:");
    #10 assign a = 64'h0230000000000000; assign b = 64'h3A80000000000000;
    #10 assign a = 64'h023FFFFFFFFFFFFF; assign b = 64'h3A8FFFFFFFFFFFFF;

    #10 $display("\n2**-987 * 2**-88:");
    #10 assign a = 64'h0240000000000000; assign b = 64'h3A70000000000000;
    #10 assign a = 64'h024FFFFFFFFFFFFF; assign b = 64'h3A7FFFFFFFFFFFFF;

    #10 $display("\n2**-986 * 2**-89:");
    #10 assign a = 64'h0250000000000000; assign b = 64'h3A60000000000000;
    #10 assign a = 64'h025FFFFFFFFFFFFF; assign b = 64'h3A6FFFFFFFFFFFFF;

    #10 $display("\n2**-985 * 2**-90:");
    #10 assign a = 64'h0260000000000000; assign b = 64'h3A50000000000000;
    #10 assign a = 64'h026FFFFFFFFFFFFF; assign b = 64'h3A5FFFFFFFFFFFFF;

    #10 $display("\n2**-984 * 2**-91:");
    #10 assign a = 64'h0270000000000000; assign b = 64'h3A40000000000000;
    #10 assign a = 64'h027FFFFFFFFFFFFF; assign b = 64'h3A4FFFFFFFFFFFFF;

    #10 $display("\n2**-983 * 2**-92:");
    #10 assign a = 64'h0280000000000000; assign b = 64'h3A30000000000000;
    #10 assign a = 64'h028FFFFFFFFFFFFF; assign b = 64'h3A3FFFFFFFFFFFFF;

    #10 $display("\n2**-982 * 2**-93:");
    #10 assign a = 64'h0290000000000000; assign b = 64'h3A20000000000000;
    #10 assign a = 64'h029FFFFFFFFFFFFF; assign b = 64'h3A2FFFFFFFFFFFFF;

    #10 $display("\n2**-981 * 2**-94:");
    #10 assign a = 64'h02A0000000000000; assign b = 64'h3A10000000000000;
    #10 assign a = 64'h02AFFFFFFFFFFFFF; assign b = 64'h3A1FFFFFFFFFFFFF;

    #10 $display("\n2**-980 * 2**-95:");
    #10 assign a = 64'h02B0000000000000; assign b = 64'h3A00000000000000;
    #10 assign a = 64'h02BFFFFFFFFFFFFF; assign b = 64'h3A0FFFFFFFFFFFFF;

    #10 $display("\n2**-979 * 2**-96:");
    #10 assign a = 64'h02C0000000000000; assign b = 64'h39F0000000000000;
    #10 assign a = 64'h02CFFFFFFFFFFFFF; assign b = 64'h39FFFFFFFFFFFFFF;

    #10 $display("\n2**-978 * 2**-97:");
    #10 assign a = 64'h02D0000000000000; assign b = 64'h39E0000000000000;
    #10 assign a = 64'h02DFFFFFFFFFFFFF; assign b = 64'h39EFFFFFFFFFFFFF;

    #10 $display("\n2**-977 * 2**-98:");
    #10 assign a = 64'h02E0000000000000; assign b = 64'h39D0000000000000;
    #10 assign a = 64'h02EFFFFFFFFFFFFF; assign b = 64'h39DFFFFFFFFFFFFF;

    #10 $display("\n2**-976 * 2**-99:");
    #10 assign a = 64'h02F0000000000000; assign b = 64'h39C0000000000000;
    #10 assign a = 64'h02FFFFFFFFFFFFFF; assign b = 64'h39CFFFFFFFFFFFFF;

    #10 $display("\n2**-975 * 2**-100:");
    #10 assign a = 64'h0300000000000000; assign b = 64'h39B0000000000000;
    #10 assign a = 64'h030FFFFFFFFFFFFF; assign b = 64'h39BFFFFFFFFFFFFF;

    #10 $display("\n2**-974 * 2**-101:");
    #10 assign a = 64'h0310000000000000; assign b = 64'h39A0000000000000;
    #10 assign a = 64'h031FFFFFFFFFFFFF; assign b = 64'h39AFFFFFFFFFFFFF;

    #10 $display("\n2**-973 * 2**-102:");
    #10 assign a = 64'h0320000000000000; assign b = 64'h3990000000000000;
    #10 assign a = 64'h032FFFFFFFFFFFFF; assign b = 64'h399FFFFFFFFFFFFF;

    #10 $display("\n2**-972 * 2**-103:");
    #10 assign a = 64'h0330000000000000; assign b = 64'h3980000000000000;
    #10 assign a = 64'h033FFFFFFFFFFFFF; assign b = 64'h398FFFFFFFFFFFFF;

    #10 $display("\n2**-971 * 2**-104:");
    #10 assign a = 64'h0340000000000000; assign b = 64'h3970000000000000;
    #10 assign a = 64'h034FFFFFFFFFFFFF; assign b = 64'h397FFFFFFFFFFFFF;

    #10 $display("\n2**-970 * 2**-105:");
    #10 assign a = 64'h0350000000000000; assign b = 64'h3960000000000000;
    #10 assign a = 64'h035FFFFFFFFFFFFF; assign b = 64'h396FFFFFFFFFFFFF;

    #10 $display("\n2**-969 * 2**-106:");
    #10 assign a = 64'h0360000000000000; assign b = 64'h3950000000000000;
    #10 assign a = 64'h036FFFFFFFFFFFFF; assign b = 64'h395FFFFFFFFFFFFF;

    #10 $display("\n2**-968 * 2**-107:");
    #10 assign a = 64'h0370000000000000; assign b = 64'h3940000000000000;
    #10 assign a = 64'h037FFFFFFFFFFFFF; assign b = 64'h394FFFFFFFFFFFFF;

    #10 $display("\n2**-967 * 2**-108:");
    #10 assign a = 64'h0380000000000000; assign b = 64'h3930000000000000;
    #10 assign a = 64'h038FFFFFFFFFFFFF; assign b = 64'h393FFFFFFFFFFFFF;

    #10 $display("\n2**-966 * 2**-109:");
    #10 assign a = 64'h0390000000000000; assign b = 64'h3920000000000000;
    #10 assign a = 64'h039FFFFFFFFFFFFF; assign b = 64'h392FFFFFFFFFFFFF;

    #10 $display("\n2**-965 * 2**-110:");
    #10 assign a = 64'h03A0000000000000; assign b = 64'h3910000000000000;
    #10 assign a = 64'h03AFFFFFFFFFFFFF; assign b = 64'h391FFFFFFFFFFFFF;

    #10 $display("\n2**-964 * 2**-111:");
    #10 assign a = 64'h03B0000000000000; assign b = 64'h3900000000000000;
    #10 assign a = 64'h03BFFFFFFFFFFFFF; assign b = 64'h390FFFFFFFFFFFFF;

    #10 $display("\n2**-963 * 2**-112:");
    #10 assign a = 64'h03C0000000000000; assign b = 64'h38F0000000000000;
    #10 assign a = 64'h03CFFFFFFFFFFFFF; assign b = 64'h38FFFFFFFFFFFFFF;

    #10 $display("\n2**-962 * 2**-113:");
    #10 assign a = 64'h03D0000000000000; assign b = 64'h38E0000000000000;
    #10 assign a = 64'h03DFFFFFFFFFFFFF; assign b = 64'h38EFFFFFFFFFFFFF;

    #10 $display("\n2**-961 * 2**-114:");
    #10 assign a = 64'h03E0000000000000; assign b = 64'h38D0000000000000;
    #10 assign a = 64'h03EFFFFFFFFFFFFF; assign b = 64'h38DFFFFFFFFFFFFF;

    #10 $display("\n2**-960 * 2**-115:");
    #10 assign a = 64'h03F0000000000000; assign b = 64'h38C0000000000000;
    #10 assign a = 64'h03FFFFFFFFFFFFFF; assign b = 64'h38CFFFFFFFFFFFFF;

    #10 $display("\n2**-959 * 2**-116:");
    #10 assign a = 64'h0400000000000000; assign b = 64'h38B0000000000000;
    #10 assign a = 64'h040FFFFFFFFFFFFF; assign b = 64'h38BFFFFFFFFFFFFF;

    #10 $display("\n2**-958 * 2**-117:");
    #10 assign a = 64'h0410000000000000; assign b = 64'h38A0000000000000;
    #10 assign a = 64'h041FFFFFFFFFFFFF; assign b = 64'h38AFFFFFFFFFFFFF;

    #10 $display("\n2**-957 * 2**-118:");
    #10 assign a = 64'h0420000000000000; assign b = 64'h3890000000000000;
    #10 assign a = 64'h042FFFFFFFFFFFFF; assign b = 64'h389FFFFFFFFFFFFF;

    #10 $display("\n2**-956 * 2**-119:");
    #10 assign a = 64'h0430000000000000; assign b = 64'h3880000000000000;
    #10 assign a = 64'h043FFFFFFFFFFFFF; assign b = 64'h388FFFFFFFFFFFFF;

    #10 $display("\n2**-955 * 2**-120:");
    #10 assign a = 64'h0440000000000000; assign b = 64'h3870000000000000;
    #10 assign a = 64'h044FFFFFFFFFFFFF; assign b = 64'h387FFFFFFFFFFFFF;

    #10 $display("\n2**-954 * 2**-121:");
    #10 assign a = 64'h0450000000000000; assign b = 64'h3860000000000000;
    #10 assign a = 64'h045FFFFFFFFFFFFF; assign b = 64'h386FFFFFFFFFFFFF;

    #10 $display("\n2**-953 * 2**-122:");
    #10 assign a = 64'h0460000000000000; assign b = 64'h3850000000000000;
    #10 assign a = 64'h046FFFFFFFFFFFFF; assign b = 64'h385FFFFFFFFFFFFF;

    #10 $display("\n2**-952 * 2**-123:");
    #10 assign a = 64'h0470000000000000; assign b = 64'h3840000000000000;
    #10 assign a = 64'h047FFFFFFFFFFFFF; assign b = 64'h384FFFFFFFFFFFFF;

    #10 $display("\n2**-951 * 2**-124:");
    #10 assign a = 64'h0480000000000000; assign b = 64'h3830000000000000;
    #10 assign a = 64'h048FFFFFFFFFFFFF; assign b = 64'h383FFFFFFFFFFFFF;

    #10 $display("\n2**-950 * 2**-125:");
    #10 assign a = 64'h0490000000000000; assign b = 64'h3820000000000000;
    #10 assign a = 64'h049FFFFFFFFFFFFF; assign b = 64'h382FFFFFFFFFFFFF;

    #10 $display("\n2**-949 * 2**-126:");
    #10 assign a = 64'h04A0000000000000; assign b = 64'h3810000000000000;
    #10 assign a = 64'h04AFFFFFFFFFFFFF; assign b = 64'h381FFFFFFFFFFFFF;

    #10 $display("\n2**-948 * 2**-127:");
    #10 assign a = 64'h04B0000000000000; assign b = 64'h3800000000000000;
    #10 assign a = 64'h04BFFFFFFFFFFFFF; assign b = 64'h380FFFFFFFFFFFFF;

    #10 $display("\n2**-947 * 2**-128:");
    #10 assign a = 64'h04C0000000000000; assign b = 64'h37F0000000000000;
    #10 assign a = 64'h04CFFFFFFFFFFFFF; assign b = 64'h37FFFFFFFFFFFFFF;

    #10 $display("\n2**-946 * 2**-129:");
    #10 assign a = 64'h04D0000000000000; assign b = 64'h37E0000000000000;
    #10 assign a = 64'h04DFFFFFFFFFFFFF; assign b = 64'h37EFFFFFFFFFFFFF;

    #10 $display("\n2**-945 * 2**-130:");
    #10 assign a = 64'h04E0000000000000; assign b = 64'h37D0000000000000;
    #10 assign a = 64'h04EFFFFFFFFFFFFF; assign b = 64'h37DFFFFFFFFFFFFF;

    #10 $display("\n2**-944 * 2**-131:");
    #10 assign a = 64'h04F0000000000000; assign b = 64'h37C0000000000000;
    #10 assign a = 64'h04FFFFFFFFFFFFFF; assign b = 64'h37CFFFFFFFFFFFFF;

    #10 $display("\n2**-943 * 2**-132:");
    #10 assign a = 64'h0500000000000000; assign b = 64'h37B0000000000000;
    #10 assign a = 64'h050FFFFFFFFFFFFF; assign b = 64'h37BFFFFFFFFFFFFF;

    #10 $display("\n2**-942 * 2**-133:");
    #10 assign a = 64'h0510000000000000; assign b = 64'h37A0000000000000;
    #10 assign a = 64'h051FFFFFFFFFFFFF; assign b = 64'h37AFFFFFFFFFFFFF;

    #10 $display("\n2**-941 * 2**-134:");
    #10 assign a = 64'h0520000000000000; assign b = 64'h3790000000000000;
    #10 assign a = 64'h052FFFFFFFFFFFFF; assign b = 64'h379FFFFFFFFFFFFF;

    #10 $display("\n2**-940 * 2**-135:");
    #10 assign a = 64'h0530000000000000; assign b = 64'h3780000000000000;
    #10 assign a = 64'h053FFFFFFFFFFFFF; assign b = 64'h378FFFFFFFFFFFFF;

    #10 $display("\n2**-939 * 2**-136:");
    #10 assign a = 64'h0540000000000000; assign b = 64'h3770000000000000;
    #10 assign a = 64'h054FFFFFFFFFFFFF; assign b = 64'h377FFFFFFFFFFFFF;

    #10 $display("\n2**-938 * 2**-137:");
    #10 assign a = 64'h0550000000000000; assign b = 64'h3760000000000000;
    #10 assign a = 64'h055FFFFFFFFFFFFF; assign b = 64'h376FFFFFFFFFFFFF;

    #10 $display("\n2**-937 * 2**-138:");
    #10 assign a = 64'h0560000000000000; assign b = 64'h3750000000000000;
    #10 assign a = 64'h056FFFFFFFFFFFFF; assign b = 64'h375FFFFFFFFFFFFF;

    #10 $display("\n2**-936 * 2**-139:");
    #10 assign a = 64'h0570000000000000; assign b = 64'h3740000000000000;
    #10 assign a = 64'h057FFFFFFFFFFFFF; assign b = 64'h374FFFFFFFFFFFFF;

    #10 $display("\n2**-935 * 2**-140:");
    #10 assign a = 64'h0580000000000000; assign b = 64'h3730000000000000;
    #10 assign a = 64'h058FFFFFFFFFFFFF; assign b = 64'h373FFFFFFFFFFFFF;

    #10 $display("\n2**-934 * 2**-141:");
    #10 assign a = 64'h0590000000000000; assign b = 64'h3720000000000000;
    #10 assign a = 64'h059FFFFFFFFFFFFF; assign b = 64'h372FFFFFFFFFFFFF;

    #10 $display("\n2**-933 * 2**-142:");
    #10 assign a = 64'h05A0000000000000; assign b = 64'h3710000000000000;
    #10 assign a = 64'h05AFFFFFFFFFFFFF; assign b = 64'h371FFFFFFFFFFFFF;

    #10 $display("\n2**-932 * 2**-143:");
    #10 assign a = 64'h05B0000000000000; assign b = 64'h3700000000000000;
    #10 assign a = 64'h05BFFFFFFFFFFFFF; assign b = 64'h370FFFFFFFFFFFFF;

    #10 $display("\n2**-931 * 2**-144:");
    #10 assign a = 64'h05C0000000000000; assign b = 64'h36F0000000000000;
    #10 assign a = 64'h05CFFFFFFFFFFFFF; assign b = 64'h36FFFFFFFFFFFFFF;

    #10 $display("\n2**-930 * 2**-145:");
    #10 assign a = 64'h05D0000000000000; assign b = 64'h36E0000000000000;
    #10 assign a = 64'h05DFFFFFFFFFFFFF; assign b = 64'h36EFFFFFFFFFFFFF;

    #10 $display("\n2**-929 * 2**-146:");
    #10 assign a = 64'h05E0000000000000; assign b = 64'h36D0000000000000;
    #10 assign a = 64'h05EFFFFFFFFFFFFF; assign b = 64'h36DFFFFFFFFFFFFF;

    #10 $display("\n2**-928 * 2**-147:");
    #10 assign a = 64'h05F0000000000000; assign b = 64'h36C0000000000000;
    #10 assign a = 64'h05FFFFFFFFFFFFFF; assign b = 64'h36CFFFFFFFFFFFFF;

    #10 $display("\n2**-927 * 2**-148:");
    #10 assign a = 64'h0600000000000000; assign b = 64'h36B0000000000000;
    #10 assign a = 64'h060FFFFFFFFFFFFF; assign b = 64'h36BFFFFFFFFFFFFF;

    #10 $display("\n2**-926 * 2**-149:");
    #10 assign a = 64'h0610000000000000; assign b = 64'h36A0000000000000;
    #10 assign a = 64'h061FFFFFFFFFFFFF; assign b = 64'h36AFFFFFFFFFFFFF;

    #10 $display("\n2**-925 * 2**-150:");
    #10 assign a = 64'h0620000000000000; assign b = 64'h3690000000000000;
    #10 assign a = 64'h062FFFFFFFFFFFFF; assign b = 64'h369FFFFFFFFFFFFF;

    #10 $display("\n2**-924 * 2**-151:");
    #10 assign a = 64'h0630000000000000; assign b = 64'h3680000000000000;
    #10 assign a = 64'h063FFFFFFFFFFFFF; assign b = 64'h368FFFFFFFFFFFFF;

    #10 $display("\n2**-923 * 2**-152:");
    #10 assign a = 64'h0640000000000000; assign b = 64'h3670000000000000;
    #10 assign a = 64'h064FFFFFFFFFFFFF; assign b = 64'h367FFFFFFFFFFFFF;

    #10 $display("\n2**-922 * 2**-153:");
    #10 assign a = 64'h0650000000000000; assign b = 64'h3660000000000000;
    #10 assign a = 64'h065FFFFFFFFFFFFF; assign b = 64'h366FFFFFFFFFFFFF;

    #10 $display("\n2**-921 * 2**-154:");
    #10 assign a = 64'h0660000000000000; assign b = 64'h3650000000000000;
    #10 assign a = 64'h066FFFFFFFFFFFFF; assign b = 64'h365FFFFFFFFFFFFF;

    #10 $display("\n2**-920 * 2**-155:");
    #10 assign a = 64'h0670000000000000; assign b = 64'h3640000000000000;
    #10 assign a = 64'h067FFFFFFFFFFFFF; assign b = 64'h364FFFFFFFFFFFFF;

    #10 $display("\n2**-919 * 2**-156:");
    #10 assign a = 64'h0680000000000000; assign b = 64'h3630000000000000;
    #10 assign a = 64'h068FFFFFFFFFFFFF; assign b = 64'h363FFFFFFFFFFFFF;

    #10 $display("\n2**-918 * 2**-157:");
    #10 assign a = 64'h0690000000000000; assign b = 64'h3620000000000000;
    #10 assign a = 64'h069FFFFFFFFFFFFF; assign b = 64'h362FFFFFFFFFFFFF;

    #10 $display("\n2**-917 * 2**-158:");
    #10 assign a = 64'h06A0000000000000; assign b = 64'h3610000000000000;
    #10 assign a = 64'h06AFFFFFFFFFFFFF; assign b = 64'h361FFFFFFFFFFFFF;

    #10 $display("\n2**-916 * 2**-159:");
    #10 assign a = 64'h06B0000000000000; assign b = 64'h3600000000000000;
    #10 assign a = 64'h06BFFFFFFFFFFFFF; assign b = 64'h360FFFFFFFFFFFFF;

    #10 $display("\n2**-915 * 2**-160:");
    #10 assign a = 64'h06C0000000000000; assign b = 64'h35F0000000000000;
    #10 assign a = 64'h06CFFFFFFFFFFFFF; assign b = 64'h35FFFFFFFFFFFFFF;

    #10 $display("\n2**-914 * 2**-161:");
    #10 assign a = 64'h06D0000000000000; assign b = 64'h35E0000000000000;
    #10 assign a = 64'h06DFFFFFFFFFFFFF; assign b = 64'h35EFFFFFFFFFFFFF;

    #10 $display("\n2**-913 * 2**-162:");
    #10 assign a = 64'h06E0000000000000; assign b = 64'h35D0000000000000;
    #10 assign a = 64'h06EFFFFFFFFFFFFF; assign b = 64'h35DFFFFFFFFFFFFF;

    #10 $display("\n2**-912 * 2**-163:");
    #10 assign a = 64'h06F0000000000000; assign b = 64'h35C0000000000000;
    #10 assign a = 64'h06FFFFFFFFFFFFFF; assign b = 64'h35CFFFFFFFFFFFFF;

    #10 $display("\n2**-911 * 2**-164:");
    #10 assign a = 64'h0700000000000000; assign b = 64'h35B0000000000000;
    #10 assign a = 64'h070FFFFFFFFFFFFF; assign b = 64'h35BFFFFFFFFFFFFF;

    #10 $display("\n2**-910 * 2**-165:");
    #10 assign a = 64'h0710000000000000; assign b = 64'h35A0000000000000;
    #10 assign a = 64'h071FFFFFFFFFFFFF; assign b = 64'h35AFFFFFFFFFFFFF;

    #10 $display("\n2**-909 * 2**-166:");
    #10 assign a = 64'h0720000000000000; assign b = 64'h3590000000000000;
    #10 assign a = 64'h072FFFFFFFFFFFFF; assign b = 64'h359FFFFFFFFFFFFF;

    #10 $display("\n2**-908 * 2**-167:");
    #10 assign a = 64'h0730000000000000; assign b = 64'h3580000000000000;
    #10 assign a = 64'h073FFFFFFFFFFFFF; assign b = 64'h358FFFFFFFFFFFFF;

    #10 $display("\n2**-907 * 2**-168:");
    #10 assign a = 64'h0740000000000000; assign b = 64'h3570000000000000;
    #10 assign a = 64'h074FFFFFFFFFFFFF; assign b = 64'h357FFFFFFFFFFFFF;

    #10 $display("\n2**-906 * 2**-169:");
    #10 assign a = 64'h0750000000000000; assign b = 64'h3560000000000000;
    #10 assign a = 64'h075FFFFFFFFFFFFF; assign b = 64'h356FFFFFFFFFFFFF;

    #10 $display("\n2**-905 * 2**-170:");
    #10 assign a = 64'h0760000000000000; assign b = 64'h3550000000000000;
    #10 assign a = 64'h076FFFFFFFFFFFFF; assign b = 64'h355FFFFFFFFFFFFF;

    #10 $display("\n2**-904 * 2**-171:");
    #10 assign a = 64'h0770000000000000; assign b = 64'h3540000000000000;
    #10 assign a = 64'h077FFFFFFFFFFFFF; assign b = 64'h354FFFFFFFFFFFFF;

    #10 $display("\n2**-903 * 2**-172:");
    #10 assign a = 64'h0780000000000000; assign b = 64'h3530000000000000;
    #10 assign a = 64'h078FFFFFFFFFFFFF; assign b = 64'h353FFFFFFFFFFFFF;

    #10 $display("\n2**-902 * 2**-173:");
    #10 assign a = 64'h0790000000000000; assign b = 64'h3520000000000000;
    #10 assign a = 64'h079FFFFFFFFFFFFF; assign b = 64'h352FFFFFFFFFFFFF;

    #10 $display("\n2**-901 * 2**-174:");
    #10 assign a = 64'h07A0000000000000; assign b = 64'h3510000000000000;
    #10 assign a = 64'h07AFFFFFFFFFFFFF; assign b = 64'h351FFFFFFFFFFFFF;

    #10 $display("\n2**-900 * 2**-175:");
    #10 assign a = 64'h07B0000000000000; assign b = 64'h3500000000000000;
    #10 assign a = 64'h07BFFFFFFFFFFFFF; assign b = 64'h350FFFFFFFFFFFFF;

    #10 $display("\n2**-899 * 2**-176:");
    #10 assign a = 64'h07C0000000000000; assign b = 64'h34F0000000000000;
    #10 assign a = 64'h07CFFFFFFFFFFFFF; assign b = 64'h34FFFFFFFFFFFFFF;

    #10 $display("\n2**-898 * 2**-177:");
    #10 assign a = 64'h07D0000000000000; assign b = 64'h34E0000000000000;
    #10 assign a = 64'h07DFFFFFFFFFFFFF; assign b = 64'h34EFFFFFFFFFFFFF;

    #10 $display("\n2**-897 * 2**-178:");
    #10 assign a = 64'h07E0000000000000; assign b = 64'h34D0000000000000;
    #10 assign a = 64'h07EFFFFFFFFFFFFF; assign b = 64'h34DFFFFFFFFFFFFF;

    #10 $display("\n2**-896 * 2**-179:");
    #10 assign a = 64'h07F0000000000000; assign b = 64'h34C0000000000000;
    #10 assign a = 64'h07FFFFFFFFFFFFFF; assign b = 64'h34CFFFFFFFFFFFFF;

    #10 $display("\n2**-895 * 2**-180:");
    #10 assign a = 64'h0800000000000000; assign b = 64'h34B0000000000000;
    #10 assign a = 64'h080FFFFFFFFFFFFF; assign b = 64'h34BFFFFFFFFFFFFF;

    #10 $display("\n2**-894 * 2**-181:");
    #10 assign a = 64'h0810000000000000; assign b = 64'h34A0000000000000;
    #10 assign a = 64'h081FFFFFFFFFFFFF; assign b = 64'h34AFFFFFFFFFFFFF;

    #10 $display("\n2**-893 * 2**-182:");
    #10 assign a = 64'h0820000000000000; assign b = 64'h3490000000000000;
    #10 assign a = 64'h082FFFFFFFFFFFFF; assign b = 64'h349FFFFFFFFFFFFF;

    #10 $display("\n2**-892 * 2**-183:");
    #10 assign a = 64'h0830000000000000; assign b = 64'h3480000000000000;
    #10 assign a = 64'h083FFFFFFFFFFFFF; assign b = 64'h348FFFFFFFFFFFFF;

    #10 $display("\n2**-891 * 2**-184:");
    #10 assign a = 64'h0840000000000000; assign b = 64'h3470000000000000;
    #10 assign a = 64'h084FFFFFFFFFFFFF; assign b = 64'h347FFFFFFFFFFFFF;

    #10 $display("\n2**-890 * 2**-185:");
    #10 assign a = 64'h0850000000000000; assign b = 64'h3460000000000000;
    #10 assign a = 64'h085FFFFFFFFFFFFF; assign b = 64'h346FFFFFFFFFFFFF;

    #10 $display("\n2**-889 * 2**-186:");
    #10 assign a = 64'h0860000000000000; assign b = 64'h3450000000000000;
    #10 assign a = 64'h086FFFFFFFFFFFFF; assign b = 64'h345FFFFFFFFFFFFF;

    #10 $display("\n2**-888 * 2**-187:");
    #10 assign a = 64'h0870000000000000; assign b = 64'h3440000000000000;
    #10 assign a = 64'h087FFFFFFFFFFFFF; assign b = 64'h344FFFFFFFFFFFFF;

    #10 $display("\n2**-887 * 2**-188:");
    #10 assign a = 64'h0880000000000000; assign b = 64'h3430000000000000;
    #10 assign a = 64'h088FFFFFFFFFFFFF; assign b = 64'h343FFFFFFFFFFFFF;

    #10 $display("\n2**-886 * 2**-189:");
    #10 assign a = 64'h0890000000000000; assign b = 64'h3420000000000000;
    #10 assign a = 64'h089FFFFFFFFFFFFF; assign b = 64'h342FFFFFFFFFFFFF;

    #10 $display("\n2**-885 * 2**-190:");
    #10 assign a = 64'h08A0000000000000; assign b = 64'h3410000000000000;
    #10 assign a = 64'h08AFFFFFFFFFFFFF; assign b = 64'h341FFFFFFFFFFFFF;

    #10 $display("\n2**-884 * 2**-191:");
    #10 assign a = 64'h08B0000000000000; assign b = 64'h3400000000000000;
    #10 assign a = 64'h08BFFFFFFFFFFFFF; assign b = 64'h340FFFFFFFFFFFFF;

    #10 $display("\n2**-883 * 2**-192:");
    #10 assign a = 64'h08C0000000000000; assign b = 64'h33F0000000000000;
    #10 assign a = 64'h08CFFFFFFFFFFFFF; assign b = 64'h33FFFFFFFFFFFFFF;

    #10 $display("\n2**-882 * 2**-193:");
    #10 assign a = 64'h08D0000000000000; assign b = 64'h33E0000000000000;
    #10 assign a = 64'h08DFFFFFFFFFFFFF; assign b = 64'h33EFFFFFFFFFFFFF;

    #10 $display("\n2**-881 * 2**-194:");
    #10 assign a = 64'h08E0000000000000; assign b = 64'h33D0000000000000;
    #10 assign a = 64'h08EFFFFFFFFFFFFF; assign b = 64'h33DFFFFFFFFFFFFF;

    #10 $display("\n2**-880 * 2**-195:");
    #10 assign a = 64'h08F0000000000000; assign b = 64'h33C0000000000000;
    #10 assign a = 64'h08FFFFFFFFFFFFFF; assign b = 64'h33CFFFFFFFFFFFFF;

    #10 $display("\n2**-879 * 2**-196:");
    #10 assign a = 64'h0900000000000000; assign b = 64'h33B0000000000000;
    #10 assign a = 64'h090FFFFFFFFFFFFF; assign b = 64'h33BFFFFFFFFFFFFF;

    #10 $display("\n2**-878 * 2**-197:");
    #10 assign a = 64'h0910000000000000; assign b = 64'h33A0000000000000;
    #10 assign a = 64'h091FFFFFFFFFFFFF; assign b = 64'h33AFFFFFFFFFFFFF;

    #10 $display("\n2**-877 * 2**-198:");
    #10 assign a = 64'h0920000000000000; assign b = 64'h3390000000000000;
    #10 assign a = 64'h092FFFFFFFFFFFFF; assign b = 64'h339FFFFFFFFFFFFF;

    #10 $display("\n2**-876 * 2**-199:");
    #10 assign a = 64'h0930000000000000; assign b = 64'h3380000000000000;
    #10 assign a = 64'h093FFFFFFFFFFFFF; assign b = 64'h338FFFFFFFFFFFFF;

    #10 $display("\n2**-875 * 2**-200:");
    #10 assign a = 64'h0940000000000000; assign b = 64'h3370000000000000;
    #10 assign a = 64'h094FFFFFFFFFFFFF; assign b = 64'h337FFFFFFFFFFFFF;

    #10 $display("\n2**-874 * 2**-201:");
    #10 assign a = 64'h0950000000000000; assign b = 64'h3360000000000000;
    #10 assign a = 64'h095FFFFFFFFFFFFF; assign b = 64'h336FFFFFFFFFFFFF;

    #10 $display("\n2**-873 * 2**-202:");
    #10 assign a = 64'h0960000000000000; assign b = 64'h3350000000000000;
    #10 assign a = 64'h096FFFFFFFFFFFFF; assign b = 64'h335FFFFFFFFFFFFF;

    #10 $display("\n2**-872 * 2**-203:");
    #10 assign a = 64'h0970000000000000; assign b = 64'h3340000000000000;
    #10 assign a = 64'h097FFFFFFFFFFFFF; assign b = 64'h334FFFFFFFFFFFFF;

    #10 $display("\n2**-871 * 2**-204:");
    #10 assign a = 64'h0980000000000000; assign b = 64'h3330000000000000;
    #10 assign a = 64'h098FFFFFFFFFFFFF; assign b = 64'h333FFFFFFFFFFFFF;

    #10 $display("\n2**-870 * 2**-205:");
    #10 assign a = 64'h0990000000000000; assign b = 64'h3320000000000000;
    #10 assign a = 64'h099FFFFFFFFFFFFF; assign b = 64'h332FFFFFFFFFFFFF;

    #10 $display("\n2**-869 * 2**-206:");
    #10 assign a = 64'h09A0000000000000; assign b = 64'h3310000000000000;
    #10 assign a = 64'h09AFFFFFFFFFFFFF; assign b = 64'h331FFFFFFFFFFFFF;

    #10 $display("\n2**-868 * 2**-207:");
    #10 assign a = 64'h09B0000000000000; assign b = 64'h3300000000000000;
    #10 assign a = 64'h09BFFFFFFFFFFFFF; assign b = 64'h330FFFFFFFFFFFFF;

    #10 $display("\n2**-867 * 2**-208:");
    #10 assign a = 64'h09C0000000000000; assign b = 64'h32F0000000000000;
    #10 assign a = 64'h09CFFFFFFFFFFFFF; assign b = 64'h32FFFFFFFFFFFFFF;

    #10 $display("\n2**-866 * 2**-209:");
    #10 assign a = 64'h09D0000000000000; assign b = 64'h32E0000000000000;
    #10 assign a = 64'h09DFFFFFFFFFFFFF; assign b = 64'h32EFFFFFFFFFFFFF;

    #10 $display("\n2**-865 * 2**-210:");
    #10 assign a = 64'h09E0000000000000; assign b = 64'h32D0000000000000;
    #10 assign a = 64'h09EFFFFFFFFFFFFF; assign b = 64'h32DFFFFFFFFFFFFF;

    #10 $display("\n2**-864 * 2**-211:");
    #10 assign a = 64'h09F0000000000000; assign b = 64'h32C0000000000000;
    #10 assign a = 64'h09FFFFFFFFFFFFFF; assign b = 64'h32CFFFFFFFFFFFFF;

    #10 $display("\n2**-863 * 2**-212:");
    #10 assign a = 64'h0A00000000000000; assign b = 64'h32B0000000000000;
    #10 assign a = 64'h0A0FFFFFFFFFFFFF; assign b = 64'h32BFFFFFFFFFFFFF;

    #10 $display("\n2**-862 * 2**-213:");
    #10 assign a = 64'h0A10000000000000; assign b = 64'h32A0000000000000;
    #10 assign a = 64'h0A1FFFFFFFFFFFFF; assign b = 64'h32AFFFFFFFFFFFFF;

    #10 $display("\n2**-861 * 2**-214:");
    #10 assign a = 64'h0A20000000000000; assign b = 64'h3290000000000000;
    #10 assign a = 64'h0A2FFFFFFFFFFFFF; assign b = 64'h329FFFFFFFFFFFFF;

    #10 $display("\n2**-860 * 2**-215:");
    #10 assign a = 64'h0A30000000000000; assign b = 64'h3280000000000000;
    #10 assign a = 64'h0A3FFFFFFFFFFFFF; assign b = 64'h328FFFFFFFFFFFFF;

    #10 $display("\n2**-859 * 2**-216:");
    #10 assign a = 64'h0A40000000000000; assign b = 64'h3270000000000000;
    #10 assign a = 64'h0A4FFFFFFFFFFFFF; assign b = 64'h327FFFFFFFFFFFFF;

    #10 $display("\n2**-858 * 2**-217:");
    #10 assign a = 64'h0A50000000000000; assign b = 64'h3260000000000000;
    #10 assign a = 64'h0A5FFFFFFFFFFFFF; assign b = 64'h326FFFFFFFFFFFFF;

    #10 $display("\n2**-857 * 2**-218:");
    #10 assign a = 64'h0A60000000000000; assign b = 64'h3250000000000000;
    #10 assign a = 64'h0A6FFFFFFFFFFFFF; assign b = 64'h325FFFFFFFFFFFFF;

    #10 $display("\n2**-856 * 2**-219:");
    #10 assign a = 64'h0A70000000000000; assign b = 64'h3240000000000000;
    #10 assign a = 64'h0A7FFFFFFFFFFFFF; assign b = 64'h324FFFFFFFFFFFFF;

    #10 $display("\n2**-855 * 2**-220:");
    #10 assign a = 64'h0A80000000000000; assign b = 64'h3230000000000000;
    #10 assign a = 64'h0A8FFFFFFFFFFFFF; assign b = 64'h323FFFFFFFFFFFFF;

    #10 $display("\n2**-854 * 2**-221:");
    #10 assign a = 64'h0A90000000000000; assign b = 64'h3220000000000000;
    #10 assign a = 64'h0A9FFFFFFFFFFFFF; assign b = 64'h322FFFFFFFFFFFFF;

    #10 $display("\n2**-853 * 2**-222:");
    #10 assign a = 64'h0AA0000000000000; assign b = 64'h3210000000000000;
    #10 assign a = 64'h0AAFFFFFFFFFFFFF; assign b = 64'h321FFFFFFFFFFFFF;

    #10 $display("\n2**-852 * 2**-223:");
    #10 assign a = 64'h0AB0000000000000; assign b = 64'h3200000000000000;
    #10 assign a = 64'h0ABFFFFFFFFFFFFF; assign b = 64'h320FFFFFFFFFFFFF;

    #10 $display("\n2**-851 * 2**-224:");
    #10 assign a = 64'h0AC0000000000000; assign b = 64'h31F0000000000000;
    #10 assign a = 64'h0ACFFFFFFFFFFFFF; assign b = 64'h31FFFFFFFFFFFFFF;

    #10 $display("\n2**-850 * 2**-225:");
    #10 assign a = 64'h0AD0000000000000; assign b = 64'h31E0000000000000;
    #10 assign a = 64'h0ADFFFFFFFFFFFFF; assign b = 64'h31EFFFFFFFFFFFFF;

    #10 $display("\n2**-849 * 2**-226:");
    #10 assign a = 64'h0AE0000000000000; assign b = 64'h31D0000000000000;
    #10 assign a = 64'h0AEFFFFFFFFFFFFF; assign b = 64'h31DFFFFFFFFFFFFF;

    #10 $display("\n2**-848 * 2**-227:");
    #10 assign a = 64'h0AF0000000000000; assign b = 64'h31C0000000000000;
    #10 assign a = 64'h0AFFFFFFFFFFFFFF; assign b = 64'h31CFFFFFFFFFFFFF;

    #10 $display("\n2**-847 * 2**-228:");
    #10 assign a = 64'h0B00000000000000; assign b = 64'h31B0000000000000;
    #10 assign a = 64'h0B0FFFFFFFFFFFFF; assign b = 64'h31BFFFFFFFFFFFFF;

    #10 $display("\n2**-846 * 2**-229:");
    #10 assign a = 64'h0B10000000000000; assign b = 64'h31A0000000000000;
    #10 assign a = 64'h0B1FFFFFFFFFFFFF; assign b = 64'h31AFFFFFFFFFFFFF;

    #10 $display("\n2**-845 * 2**-230:");
    #10 assign a = 64'h0B20000000000000; assign b = 64'h3190000000000000;
    #10 assign a = 64'h0B2FFFFFFFFFFFFF; assign b = 64'h319FFFFFFFFFFFFF;

    #10 $display("\n2**-844 * 2**-231:");
    #10 assign a = 64'h0B30000000000000; assign b = 64'h3180000000000000;
    #10 assign a = 64'h0B3FFFFFFFFFFFFF; assign b = 64'h318FFFFFFFFFFFFF;

    #10 $display("\n2**-843 * 2**-232:");
    #10 assign a = 64'h0B40000000000000; assign b = 64'h3170000000000000;
    #10 assign a = 64'h0B4FFFFFFFFFFFFF; assign b = 64'h317FFFFFFFFFFFFF;

    #10 $display("\n2**-842 * 2**-233:");
    #10 assign a = 64'h0B50000000000000; assign b = 64'h3160000000000000;
    #10 assign a = 64'h0B5FFFFFFFFFFFFF; assign b = 64'h316FFFFFFFFFFFFF;

    #10 $display("\n2**-841 * 2**-234:");
    #10 assign a = 64'h0B60000000000000; assign b = 64'h3150000000000000;
    #10 assign a = 64'h0B6FFFFFFFFFFFFF; assign b = 64'h315FFFFFFFFFFFFF;

    #10 $display("\n2**-840 * 2**-235:");
    #10 assign a = 64'h0B70000000000000; assign b = 64'h3140000000000000;
    #10 assign a = 64'h0B7FFFFFFFFFFFFF; assign b = 64'h314FFFFFFFFFFFFF;

    #10 $display("\n2**-839 * 2**-236:");
    #10 assign a = 64'h0B80000000000000; assign b = 64'h3130000000000000;
    #10 assign a = 64'h0B8FFFFFFFFFFFFF; assign b = 64'h313FFFFFFFFFFFFF;

    #10 $display("\n2**-838 * 2**-237:");
    #10 assign a = 64'h0B90000000000000; assign b = 64'h3120000000000000;
    #10 assign a = 64'h0B9FFFFFFFFFFFFF; assign b = 64'h312FFFFFFFFFFFFF;

    #10 $display("\n2**-837 * 2**-238:");
    #10 assign a = 64'h0BA0000000000000; assign b = 64'h3110000000000000;
    #10 assign a = 64'h0BAFFFFFFFFFFFFF; assign b = 64'h311FFFFFFFFFFFFF;

    #10 $display("\n2**-836 * 2**-239:");
    #10 assign a = 64'h0BB0000000000000; assign b = 64'h3100000000000000;
    #10 assign a = 64'h0BBFFFFFFFFFFFFF; assign b = 64'h310FFFFFFFFFFFFF;

    #10 $display("\n2**-835 * 2**-240:");
    #10 assign a = 64'h0BC0000000000000; assign b = 64'h30F0000000000000;
    #10 assign a = 64'h0BCFFFFFFFFFFFFF; assign b = 64'h30FFFFFFFFFFFFFF;

    #10 $display("\n2**-834 * 2**-241:");
    #10 assign a = 64'h0BD0000000000000; assign b = 64'h30E0000000000000;
    #10 assign a = 64'h0BDFFFFFFFFFFFFF; assign b = 64'h30EFFFFFFFFFFFFF;

    #10 $display("\n2**-833 * 2**-242:");
    #10 assign a = 64'h0BE0000000000000; assign b = 64'h30D0000000000000;
    #10 assign a = 64'h0BEFFFFFFFFFFFFF; assign b = 64'h30DFFFFFFFFFFFFF;

    #10 $display("\n2**-832 * 2**-243:");
    #10 assign a = 64'h0BF0000000000000; assign b = 64'h30C0000000000000;
    #10 assign a = 64'h0BFFFFFFFFFFFFFF; assign b = 64'h30CFFFFFFFFFFFFF;

    #10 $display("\n2**-831 * 2**-244:");
    #10 assign a = 64'h0C00000000000000; assign b = 64'h30B0000000000000;
    #10 assign a = 64'h0C0FFFFFFFFFFFFF; assign b = 64'h30BFFFFFFFFFFFFF;

    #10 $display("\n2**-830 * 2**-245:");
    #10 assign a = 64'h0C10000000000000; assign b = 64'h30A0000000000000;
    #10 assign a = 64'h0C1FFFFFFFFFFFFF; assign b = 64'h30AFFFFFFFFFFFFF;

    #10 $display("\n2**-829 * 2**-246:");
    #10 assign a = 64'h0C20000000000000; assign b = 64'h3090000000000000;
    #10 assign a = 64'h0C2FFFFFFFFFFFFF; assign b = 64'h309FFFFFFFFFFFFF;

    #10 $display("\n2**-828 * 2**-247:");
    #10 assign a = 64'h0C30000000000000; assign b = 64'h3080000000000000;
    #10 assign a = 64'h0C3FFFFFFFFFFFFF; assign b = 64'h308FFFFFFFFFFFFF;

    #10 $display("\n2**-827 * 2**-248:");
    #10 assign a = 64'h0C40000000000000; assign b = 64'h3070000000000000;
    #10 assign a = 64'h0C4FFFFFFFFFFFFF; assign b = 64'h307FFFFFFFFFFFFF;

    #10 $display("\n2**-826 * 2**-249:");
    #10 assign a = 64'h0C50000000000000; assign b = 64'h3060000000000000;
    #10 assign a = 64'h0C5FFFFFFFFFFFFF; assign b = 64'h306FFFFFFFFFFFFF;

    #10 $display("\n2**-825 * 2**-250:");
    #10 assign a = 64'h0C60000000000000; assign b = 64'h3050000000000000;
    #10 assign a = 64'h0C6FFFFFFFFFFFFF; assign b = 64'h305FFFFFFFFFFFFF;

    #10 $display("\n2**-824 * 2**-251:");
    #10 assign a = 64'h0C70000000000000; assign b = 64'h3040000000000000;
    #10 assign a = 64'h0C7FFFFFFFFFFFFF; assign b = 64'h304FFFFFFFFFFFFF;

    #10 $display("\n2**-823 * 2**-252:");
    #10 assign a = 64'h0C80000000000000; assign b = 64'h3030000000000000;
    #10 assign a = 64'h0C8FFFFFFFFFFFFF; assign b = 64'h303FFFFFFFFFFFFF;

    #10 $display("\n2**-822 * 2**-253:");
    #10 assign a = 64'h0C90000000000000; assign b = 64'h3020000000000000;
    #10 assign a = 64'h0C9FFFFFFFFFFFFF; assign b = 64'h302FFFFFFFFFFFFF;

    #10 $display("\n2**-821 * 2**-254:");
    #10 assign a = 64'h0CA0000000000000; assign b = 64'h3010000000000000;
    #10 assign a = 64'h0CAFFFFFFFFFFFFF; assign b = 64'h301FFFFFFFFFFFFF;

    #10 $display("\n2**-820 * 2**-255:");
    #10 assign a = 64'h0CB0000000000000; assign b = 64'h3000000000000000;
    #10 assign a = 64'h0CBFFFFFFFFFFFFF; assign b = 64'h300FFFFFFFFFFFFF;

    #10 $display("\n2**-819 * 2**-256:");
    #10 assign a = 64'h0CC0000000000000; assign b = 64'h2FF0000000000000;
    #10 assign a = 64'h0CCFFFFFFFFFFFFF; assign b = 64'h2FFFFFFFFFFFFFFF;

    #10 $display("\n2**-818 * 2**-257:");
    #10 assign a = 64'h0CD0000000000000; assign b = 64'h2FE0000000000000;
    #10 assign a = 64'h0CDFFFFFFFFFFFFF; assign b = 64'h2FEFFFFFFFFFFFFF;

    #10 $display("\n2**-817 * 2**-258:");
    #10 assign a = 64'h0CE0000000000000; assign b = 64'h2FD0000000000000;
    #10 assign a = 64'h0CEFFFFFFFFFFFFF; assign b = 64'h2FDFFFFFFFFFFFFF;

    #10 $display("\n2**-816 * 2**-259:");
    #10 assign a = 64'h0CF0000000000000; assign b = 64'h2FC0000000000000;
    #10 assign a = 64'h0CFFFFFFFFFFFFFF; assign b = 64'h2FCFFFFFFFFFFFFF;

    #10 $display("\n2**-815 * 2**-260:");
    #10 assign a = 64'h0D00000000000000; assign b = 64'h2FB0000000000000;
    #10 assign a = 64'h0D0FFFFFFFFFFFFF; assign b = 64'h2FBFFFFFFFFFFFFF;

    #10 $display("\n2**-814 * 2**-261:");
    #10 assign a = 64'h0D10000000000000; assign b = 64'h2FA0000000000000;
    #10 assign a = 64'h0D1FFFFFFFFFFFFF; assign b = 64'h2FAFFFFFFFFFFFFF;

    #10 $display("\n2**-813 * 2**-262:");
    #10 assign a = 64'h0D20000000000000; assign b = 64'h2F90000000000000;
    #10 assign a = 64'h0D2FFFFFFFFFFFFF; assign b = 64'h2F9FFFFFFFFFFFFF;

    #10 $display("\n2**-812 * 2**-263:");
    #10 assign a = 64'h0D30000000000000; assign b = 64'h2F80000000000000;
    #10 assign a = 64'h0D3FFFFFFFFFFFFF; assign b = 64'h2F8FFFFFFFFFFFFF;

    #10 $display("\n2**-811 * 2**-264:");
    #10 assign a = 64'h0D40000000000000; assign b = 64'h2F70000000000000;
    #10 assign a = 64'h0D4FFFFFFFFFFFFF; assign b = 64'h2F7FFFFFFFFFFFFF;

    #10 $display("\n2**-810 * 2**-265:");
    #10 assign a = 64'h0D50000000000000; assign b = 64'h2F60000000000000;
    #10 assign a = 64'h0D5FFFFFFFFFFFFF; assign b = 64'h2F6FFFFFFFFFFFFF;

    #10 $display("\n2**-809 * 2**-266:");
    #10 assign a = 64'h0D60000000000000; assign b = 64'h2F50000000000000;
    #10 assign a = 64'h0D6FFFFFFFFFFFFF; assign b = 64'h2F5FFFFFFFFFFFFF;

    #10 $display("\n2**-808 * 2**-267:");
    #10 assign a = 64'h0D70000000000000; assign b = 64'h2F40000000000000;
    #10 assign a = 64'h0D7FFFFFFFFFFFFF; assign b = 64'h2F4FFFFFFFFFFFFF;

    #10 $display("\n2**-807 * 2**-268:");
    #10 assign a = 64'h0D80000000000000; assign b = 64'h2F30000000000000;
    #10 assign a = 64'h0D8FFFFFFFFFFFFF; assign b = 64'h2F3FFFFFFFFFFFFF;

    #10 $display("\n2**-806 * 2**-269:");
    #10 assign a = 64'h0D90000000000000; assign b = 64'h2F20000000000000;
    #10 assign a = 64'h0D9FFFFFFFFFFFFF; assign b = 64'h2F2FFFFFFFFFFFFF;

    #10 $display("\n2**-805 * 2**-270:");
    #10 assign a = 64'h0DA0000000000000; assign b = 64'h2F10000000000000;
    #10 assign a = 64'h0DAFFFFFFFFFFFFF; assign b = 64'h2F1FFFFFFFFFFFFF;

    #10 $display("\n2**-804 * 2**-271:");
    #10 assign a = 64'h0DB0000000000000; assign b = 64'h2F00000000000000;
    #10 assign a = 64'h0DBFFFFFFFFFFFFF; assign b = 64'h2F0FFFFFFFFFFFFF;

    #10 $display("\n2**-803 * 2**-272:");
    #10 assign a = 64'h0DC0000000000000; assign b = 64'h2EF0000000000000;
    #10 assign a = 64'h0DCFFFFFFFFFFFFF; assign b = 64'h2EFFFFFFFFFFFFFF;

    #10 $display("\n2**-802 * 2**-273:");
    #10 assign a = 64'h0DD0000000000000; assign b = 64'h2EE0000000000000;
    #10 assign a = 64'h0DDFFFFFFFFFFFFF; assign b = 64'h2EEFFFFFFFFFFFFF;

    #10 $display("\n2**-801 * 2**-274:");
    #10 assign a = 64'h0DE0000000000000; assign b = 64'h2ED0000000000000;
    #10 assign a = 64'h0DEFFFFFFFFFFFFF; assign b = 64'h2EDFFFFFFFFFFFFF;

    #10 $display("\n2**-800 * 2**-275:");
    #10 assign a = 64'h0DF0000000000000; assign b = 64'h2EC0000000000000;
    #10 assign a = 64'h0DFFFFFFFFFFFFFF; assign b = 64'h2ECFFFFFFFFFFFFF;

    #10 $display("\n2**-799 * 2**-276:");
    #10 assign a = 64'h0E00000000000000; assign b = 64'h2EB0000000000000;
    #10 assign a = 64'h0E0FFFFFFFFFFFFF; assign b = 64'h2EBFFFFFFFFFFFFF;

    #10 $display("\n2**-798 * 2**-277:");
    #10 assign a = 64'h0E10000000000000; assign b = 64'h2EA0000000000000;
    #10 assign a = 64'h0E1FFFFFFFFFFFFF; assign b = 64'h2EAFFFFFFFFFFFFF;

    #10 $display("\n2**-797 * 2**-278:");
    #10 assign a = 64'h0E20000000000000; assign b = 64'h2E90000000000000;
    #10 assign a = 64'h0E2FFFFFFFFFFFFF; assign b = 64'h2E9FFFFFFFFFFFFF;

    #10 $display("\n2**-796 * 2**-279:");
    #10 assign a = 64'h0E30000000000000; assign b = 64'h2E80000000000000;
    #10 assign a = 64'h0E3FFFFFFFFFFFFF; assign b = 64'h2E8FFFFFFFFFFFFF;

    #10 $display("\n2**-795 * 2**-280:");
    #10 assign a = 64'h0E40000000000000; assign b = 64'h2E70000000000000;
    #10 assign a = 64'h0E4FFFFFFFFFFFFF; assign b = 64'h2E7FFFFFFFFFFFFF;

    #10 $display("\n2**-794 * 2**-281:");
    #10 assign a = 64'h0E50000000000000; assign b = 64'h2E60000000000000;
    #10 assign a = 64'h0E5FFFFFFFFFFFFF; assign b = 64'h2E6FFFFFFFFFFFFF;

    #10 $display("\n2**-793 * 2**-282:");
    #10 assign a = 64'h0E60000000000000; assign b = 64'h2E50000000000000;
    #10 assign a = 64'h0E6FFFFFFFFFFFFF; assign b = 64'h2E5FFFFFFFFFFFFF;

    #10 $display("\n2**-792 * 2**-283:");
    #10 assign a = 64'h0E70000000000000; assign b = 64'h2E40000000000000;
    #10 assign a = 64'h0E7FFFFFFFFFFFFF; assign b = 64'h2E4FFFFFFFFFFFFF;

    #10 $display("\n2**-791 * 2**-284:");
    #10 assign a = 64'h0E80000000000000; assign b = 64'h2E30000000000000;
    #10 assign a = 64'h0E8FFFFFFFFFFFFF; assign b = 64'h2E3FFFFFFFFFFFFF;

    #10 $display("\n2**-790 * 2**-285:");
    #10 assign a = 64'h0E90000000000000; assign b = 64'h2E20000000000000;
    #10 assign a = 64'h0E9FFFFFFFFFFFFF; assign b = 64'h2E2FFFFFFFFFFFFF;

    #10 $display("\n2**-789 * 2**-286:");
    #10 assign a = 64'h0EA0000000000000; assign b = 64'h2E10000000000000;
    #10 assign a = 64'h0EAFFFFFFFFFFFFF; assign b = 64'h2E1FFFFFFFFFFFFF;

    #10 $display("\n2**-788 * 2**-287:");
    #10 assign a = 64'h0EB0000000000000; assign b = 64'h2E00000000000000;
    #10 assign a = 64'h0EBFFFFFFFFFFFFF; assign b = 64'h2E0FFFFFFFFFFFFF;

    #10 $display("\n2**-787 * 2**-288:");
    #10 assign a = 64'h0EC0000000000000; assign b = 64'h2DF0000000000000;
    #10 assign a = 64'h0ECFFFFFFFFFFFFF; assign b = 64'h2DFFFFFFFFFFFFFF;

    #10 $display("\n2**-786 * 2**-289:");
    #10 assign a = 64'h0ED0000000000000; assign b = 64'h2DE0000000000000;
    #10 assign a = 64'h0EDFFFFFFFFFFFFF; assign b = 64'h2DEFFFFFFFFFFFFF;

    #10 $display("\n2**-785 * 2**-290:");
    #10 assign a = 64'h0EE0000000000000; assign b = 64'h2DD0000000000000;
    #10 assign a = 64'h0EEFFFFFFFFFFFFF; assign b = 64'h2DDFFFFFFFFFFFFF;

    #10 $display("\n2**-784 * 2**-291:");
    #10 assign a = 64'h0EF0000000000000; assign b = 64'h2DC0000000000000;
    #10 assign a = 64'h0EFFFFFFFFFFFFFF; assign b = 64'h2DCFFFFFFFFFFFFF;

    #10 $display("\n2**-783 * 2**-292:");
    #10 assign a = 64'h0F00000000000000; assign b = 64'h2DB0000000000000;
    #10 assign a = 64'h0F0FFFFFFFFFFFFF; assign b = 64'h2DBFFFFFFFFFFFFF;

    #10 $display("\n2**-782 * 2**-293:");
    #10 assign a = 64'h0F10000000000000; assign b = 64'h2DA0000000000000;
    #10 assign a = 64'h0F1FFFFFFFFFFFFF; assign b = 64'h2DAFFFFFFFFFFFFF;

    #10 $display("\n2**-781 * 2**-294:");
    #10 assign a = 64'h0F20000000000000; assign b = 64'h2D90000000000000;
    #10 assign a = 64'h0F2FFFFFFFFFFFFF; assign b = 64'h2D9FFFFFFFFFFFFF;

    #10 $display("\n2**-780 * 2**-295:");
    #10 assign a = 64'h0F30000000000000; assign b = 64'h2D80000000000000;
    #10 assign a = 64'h0F3FFFFFFFFFFFFF; assign b = 64'h2D8FFFFFFFFFFFFF;

    #10 $display("\n2**-779 * 2**-296:");
    #10 assign a = 64'h0F40000000000000; assign b = 64'h2D70000000000000;
    #10 assign a = 64'h0F4FFFFFFFFFFFFF; assign b = 64'h2D7FFFFFFFFFFFFF;

    #10 $display("\n2**-778 * 2**-297:");
    #10 assign a = 64'h0F50000000000000; assign b = 64'h2D60000000000000;
    #10 assign a = 64'h0F5FFFFFFFFFFFFF; assign b = 64'h2D6FFFFFFFFFFFFF;

    #10 $display("\n2**-777 * 2**-298:");
    #10 assign a = 64'h0F60000000000000; assign b = 64'h2D50000000000000;
    #10 assign a = 64'h0F6FFFFFFFFFFFFF; assign b = 64'h2D5FFFFFFFFFFFFF;

    #10 $display("\n2**-776 * 2**-299:");
    #10 assign a = 64'h0F70000000000000; assign b = 64'h2D40000000000000;
    #10 assign a = 64'h0F7FFFFFFFFFFFFF; assign b = 64'h2D4FFFFFFFFFFFFF;

    #10 $display("\n2**-775 * 2**-300:");
    #10 assign a = 64'h0F80000000000000; assign b = 64'h2D30000000000000;
    #10 assign a = 64'h0F8FFFFFFFFFFFFF; assign b = 64'h2D3FFFFFFFFFFFFF;

    #10 $display("\n2**-774 * 2**-301:");
    #10 assign a = 64'h0F90000000000000; assign b = 64'h2D20000000000000;
    #10 assign a = 64'h0F9FFFFFFFFFFFFF; assign b = 64'h2D2FFFFFFFFFFFFF;

    #10 $display("\n2**-773 * 2**-302:");
    #10 assign a = 64'h0FA0000000000000; assign b = 64'h2D10000000000000;
    #10 assign a = 64'h0FAFFFFFFFFFFFFF; assign b = 64'h2D1FFFFFFFFFFFFF;

    #10 $display("\n2**-772 * 2**-303:");
    #10 assign a = 64'h0FB0000000000000; assign b = 64'h2D00000000000000;
    #10 assign a = 64'h0FBFFFFFFFFFFFFF; assign b = 64'h2D0FFFFFFFFFFFFF;

    #10 $display("\n2**-771 * 2**-304:");
    #10 assign a = 64'h0FC0000000000000; assign b = 64'h2CF0000000000000;
    #10 assign a = 64'h0FCFFFFFFFFFFFFF; assign b = 64'h2CFFFFFFFFFFFFFF;

    #10 $display("\n2**-770 * 2**-305:");
    #10 assign a = 64'h0FD0000000000000; assign b = 64'h2CE0000000000000;
    #10 assign a = 64'h0FDFFFFFFFFFFFFF; assign b = 64'h2CEFFFFFFFFFFFFF;

    #10 $display("\n2**-769 * 2**-306:");
    #10 assign a = 64'h0FE0000000000000; assign b = 64'h2CD0000000000000;
    #10 assign a = 64'h0FEFFFFFFFFFFFFF; assign b = 64'h2CDFFFFFFFFFFFFF;

    #10 $display("\n2**-768 * 2**-307:");
    #10 assign a = 64'h0FF0000000000000; assign b = 64'h2CC0000000000000;
    #10 assign a = 64'h0FFFFFFFFFFFFFFF; assign b = 64'h2CCFFFFFFFFFFFFF;

    #10 $display("\n2**-767 * 2**-308:");
    #10 assign a = 64'h1000000000000000; assign b = 64'h2CB0000000000000;
    #10 assign a = 64'h100FFFFFFFFFFFFF; assign b = 64'h2CBFFFFFFFFFFFFF;

    #10 $display("\n2**-766 * 2**-309:");
    #10 assign a = 64'h1010000000000000; assign b = 64'h2CA0000000000000;
    #10 assign a = 64'h101FFFFFFFFFFFFF; assign b = 64'h2CAFFFFFFFFFFFFF;

    #10 $display("\n2**-765 * 2**-310:");
    #10 assign a = 64'h1020000000000000; assign b = 64'h2C90000000000000;
    #10 assign a = 64'h102FFFFFFFFFFFFF; assign b = 64'h2C9FFFFFFFFFFFFF;

    #10 $display("\n2**-764 * 2**-311:");
    #10 assign a = 64'h1030000000000000; assign b = 64'h2C80000000000000;
    #10 assign a = 64'h103FFFFFFFFFFFFF; assign b = 64'h2C8FFFFFFFFFFFFF;

    #10 $display("\n2**-763 * 2**-312:");
    #10 assign a = 64'h1040000000000000; assign b = 64'h2C70000000000000;
    #10 assign a = 64'h104FFFFFFFFFFFFF; assign b = 64'h2C7FFFFFFFFFFFFF;

    #10 $display("\n2**-762 * 2**-313:");
    #10 assign a = 64'h1050000000000000; assign b = 64'h2C60000000000000;
    #10 assign a = 64'h105FFFFFFFFFFFFF; assign b = 64'h2C6FFFFFFFFFFFFF;

    #10 $display("\n2**-761 * 2**-314:");
    #10 assign a = 64'h1060000000000000; assign b = 64'h2C50000000000000;
    #10 assign a = 64'h106FFFFFFFFFFFFF; assign b = 64'h2C5FFFFFFFFFFFFF;

    #10 $display("\n2**-760 * 2**-315:");
    #10 assign a = 64'h1070000000000000; assign b = 64'h2C40000000000000;
    #10 assign a = 64'h107FFFFFFFFFFFFF; assign b = 64'h2C4FFFFFFFFFFFFF;

    #10 $display("\n2**-759 * 2**-316:");
    #10 assign a = 64'h1080000000000000; assign b = 64'h2C30000000000000;
    #10 assign a = 64'h108FFFFFFFFFFFFF; assign b = 64'h2C3FFFFFFFFFFFFF;

    #10 $display("\n2**-758 * 2**-317:");
    #10 assign a = 64'h1090000000000000; assign b = 64'h2C20000000000000;
    #10 assign a = 64'h109FFFFFFFFFFFFF; assign b = 64'h2C2FFFFFFFFFFFFF;

    #10 $display("\n2**-757 * 2**-318:");
    #10 assign a = 64'h10A0000000000000; assign b = 64'h2C10000000000000;
    #10 assign a = 64'h10AFFFFFFFFFFFFF; assign b = 64'h2C1FFFFFFFFFFFFF;

    #10 $display("\n2**-756 * 2**-319:");
    #10 assign a = 64'h10B0000000000000; assign b = 64'h2C00000000000000;
    #10 assign a = 64'h10BFFFFFFFFFFFFF; assign b = 64'h2C0FFFFFFFFFFFFF;

    #10 $display("\n2**-755 * 2**-320:");
    #10 assign a = 64'h10C0000000000000; assign b = 64'h2BF0000000000000;
    #10 assign a = 64'h10CFFFFFFFFFFFFF; assign b = 64'h2BFFFFFFFFFFFFFF;

    #10 $display("\n2**-754 * 2**-321:");
    #10 assign a = 64'h10D0000000000000; assign b = 64'h2BE0000000000000;
    #10 assign a = 64'h10DFFFFFFFFFFFFF; assign b = 64'h2BEFFFFFFFFFFFFF;

    #10 $display("\n2**-753 * 2**-322:");
    #10 assign a = 64'h10E0000000000000; assign b = 64'h2BD0000000000000;
    #10 assign a = 64'h10EFFFFFFFFFFFFF; assign b = 64'h2BDFFFFFFFFFFFFF;

    #10 $display("\n2**-752 * 2**-323:");
    #10 assign a = 64'h10F0000000000000; assign b = 64'h2BC0000000000000;
    #10 assign a = 64'h10FFFFFFFFFFFFFF; assign b = 64'h2BCFFFFFFFFFFFFF;

    #10 $display("\n2**-751 * 2**-324:");
    #10 assign a = 64'h1100000000000000; assign b = 64'h2BB0000000000000;
    #10 assign a = 64'h110FFFFFFFFFFFFF; assign b = 64'h2BBFFFFFFFFFFFFF;

    #10 $display("\n2**-750 * 2**-325:");
    #10 assign a = 64'h1110000000000000; assign b = 64'h2BA0000000000000;
    #10 assign a = 64'h111FFFFFFFFFFFFF; assign b = 64'h2BAFFFFFFFFFFFFF;

    #10 $display("\n2**-749 * 2**-326:");
    #10 assign a = 64'h1120000000000000; assign b = 64'h2B90000000000000;
    #10 assign a = 64'h112FFFFFFFFFFFFF; assign b = 64'h2B9FFFFFFFFFFFFF;

    #10 $display("\n2**-748 * 2**-327:");
    #10 assign a = 64'h1130000000000000; assign b = 64'h2B80000000000000;
    #10 assign a = 64'h113FFFFFFFFFFFFF; assign b = 64'h2B8FFFFFFFFFFFFF;

    #10 $display("\n2**-747 * 2**-328:");
    #10 assign a = 64'h1140000000000000; assign b = 64'h2B70000000000000;
    #10 assign a = 64'h114FFFFFFFFFFFFF; assign b = 64'h2B7FFFFFFFFFFFFF;

    #10 $display("\n2**-746 * 2**-329:");
    #10 assign a = 64'h1150000000000000; assign b = 64'h2B60000000000000;
    #10 assign a = 64'h115FFFFFFFFFFFFF; assign b = 64'h2B6FFFFFFFFFFFFF;

    #10 $display("\n2**-745 * 2**-330:");
    #10 assign a = 64'h1160000000000000; assign b = 64'h2B50000000000000;
    #10 assign a = 64'h116FFFFFFFFFFFFF; assign b = 64'h2B5FFFFFFFFFFFFF;

    #10 $display("\n2**-744 * 2**-331:");
    #10 assign a = 64'h1170000000000000; assign b = 64'h2B40000000000000;
    #10 assign a = 64'h117FFFFFFFFFFFFF; assign b = 64'h2B4FFFFFFFFFFFFF;

    #10 $display("\n2**-743 * 2**-332:");
    #10 assign a = 64'h1180000000000000; assign b = 64'h2B30000000000000;
    #10 assign a = 64'h118FFFFFFFFFFFFF; assign b = 64'h2B3FFFFFFFFFFFFF;

    #10 $display("\n2**-742 * 2**-333:");
    #10 assign a = 64'h1190000000000000; assign b = 64'h2B20000000000000;
    #10 assign a = 64'h119FFFFFFFFFFFFF; assign b = 64'h2B2FFFFFFFFFFFFF;

    #10 $display("\n2**-741 * 2**-334:");
    #10 assign a = 64'h11A0000000000000; assign b = 64'h2B10000000000000;
    #10 assign a = 64'h11AFFFFFFFFFFFFF; assign b = 64'h2B1FFFFFFFFFFFFF;

    #10 $display("\n2**-740 * 2**-335:");
    #10 assign a = 64'h11B0000000000000; assign b = 64'h2B00000000000000;
    #10 assign a = 64'h11BFFFFFFFFFFFFF; assign b = 64'h2B0FFFFFFFFFFFFF;

    #10 $display("\n2**-739 * 2**-336:");
    #10 assign a = 64'h11C0000000000000; assign b = 64'h2AF0000000000000;
    #10 assign a = 64'h11CFFFFFFFFFFFFF; assign b = 64'h2AFFFFFFFFFFFFFF;

    #10 $display("\n2**-738 * 2**-337:");
    #10 assign a = 64'h11D0000000000000; assign b = 64'h2AE0000000000000;
    #10 assign a = 64'h11DFFFFFFFFFFFFF; assign b = 64'h2AEFFFFFFFFFFFFF;

    #10 $display("\n2**-737 * 2**-338:");
    #10 assign a = 64'h11E0000000000000; assign b = 64'h2AD0000000000000;
    #10 assign a = 64'h11EFFFFFFFFFFFFF; assign b = 64'h2ADFFFFFFFFFFFFF;

    #10 $display("\n2**-736 * 2**-339:");
    #10 assign a = 64'h11F0000000000000; assign b = 64'h2AC0000000000000;
    #10 assign a = 64'h11FFFFFFFFFFFFFF; assign b = 64'h2ACFFFFFFFFFFFFF;

    #10 $display("\n2**-735 * 2**-340:");
    #10 assign a = 64'h1200000000000000; assign b = 64'h2AB0000000000000;
    #10 assign a = 64'h120FFFFFFFFFFFFF; assign b = 64'h2ABFFFFFFFFFFFFF;

    #10 $display("\n2**-734 * 2**-341:");
    #10 assign a = 64'h1210000000000000; assign b = 64'h2AA0000000000000;
    #10 assign a = 64'h121FFFFFFFFFFFFF; assign b = 64'h2AAFFFFFFFFFFFFF;

    #10 $display("\n2**-733 * 2**-342:");
    #10 assign a = 64'h1220000000000000; assign b = 64'h2A90000000000000;
    #10 assign a = 64'h122FFFFFFFFFFFFF; assign b = 64'h2A9FFFFFFFFFFFFF;

    #10 $display("\n2**-732 * 2**-343:");
    #10 assign a = 64'h1230000000000000; assign b = 64'h2A80000000000000;
    #10 assign a = 64'h123FFFFFFFFFFFFF; assign b = 64'h2A8FFFFFFFFFFFFF;

    #10 $display("\n2**-731 * 2**-344:");
    #10 assign a = 64'h1240000000000000; assign b = 64'h2A70000000000000;
    #10 assign a = 64'h124FFFFFFFFFFFFF; assign b = 64'h2A7FFFFFFFFFFFFF;

    #10 $display("\n2**-730 * 2**-345:");
    #10 assign a = 64'h1250000000000000; assign b = 64'h2A60000000000000;
    #10 assign a = 64'h125FFFFFFFFFFFFF; assign b = 64'h2A6FFFFFFFFFFFFF;

    #10 $display("\n2**-729 * 2**-346:");
    #10 assign a = 64'h1260000000000000; assign b = 64'h2A50000000000000;
    #10 assign a = 64'h126FFFFFFFFFFFFF; assign b = 64'h2A5FFFFFFFFFFFFF;

    #10 $display("\n2**-728 * 2**-347:");
    #10 assign a = 64'h1270000000000000; assign b = 64'h2A40000000000000;
    #10 assign a = 64'h127FFFFFFFFFFFFF; assign b = 64'h2A4FFFFFFFFFFFFF;

    #10 $display("\n2**-727 * 2**-348:");
    #10 assign a = 64'h1280000000000000; assign b = 64'h2A30000000000000;
    #10 assign a = 64'h128FFFFFFFFFFFFF; assign b = 64'h2A3FFFFFFFFFFFFF;

    #10 $display("\n2**-726 * 2**-349:");
    #10 assign a = 64'h1290000000000000; assign b = 64'h2A20000000000000;
    #10 assign a = 64'h129FFFFFFFFFFFFF; assign b = 64'h2A2FFFFFFFFFFFFF;

    #10 $display("\n2**-725 * 2**-350:");
    #10 assign a = 64'h12A0000000000000; assign b = 64'h2A10000000000000;
    #10 assign a = 64'h12AFFFFFFFFFFFFF; assign b = 64'h2A1FFFFFFFFFFFFF;

    #10 $display("\n2**-724 * 2**-351:");
    #10 assign a = 64'h12B0000000000000; assign b = 64'h2A00000000000000;
    #10 assign a = 64'h12BFFFFFFFFFFFFF; assign b = 64'h2A0FFFFFFFFFFFFF;

    #10 $display("\n2**-723 * 2**-352:");
    #10 assign a = 64'h12C0000000000000; assign b = 64'h29F0000000000000;
    #10 assign a = 64'h12CFFFFFFFFFFFFF; assign b = 64'h29FFFFFFFFFFFFFF;

    #10 $display("\n2**-722 * 2**-353:");
    #10 assign a = 64'h12D0000000000000; assign b = 64'h29E0000000000000;
    #10 assign a = 64'h12DFFFFFFFFFFFFF; assign b = 64'h29EFFFFFFFFFFFFF;

    #10 $display("\n2**-721 * 2**-354:");
    #10 assign a = 64'h12E0000000000000; assign b = 64'h29D0000000000000;
    #10 assign a = 64'h12EFFFFFFFFFFFFF; assign b = 64'h29DFFFFFFFFFFFFF;

    #10 $display("\n2**-720 * 2**-355:");
    #10 assign a = 64'h12F0000000000000; assign b = 64'h29C0000000000000;
    #10 assign a = 64'h12FFFFFFFFFFFFFF; assign b = 64'h29CFFFFFFFFFFFFF;

    #10 $display("\n2**-719 * 2**-356:");
    #10 assign a = 64'h1300000000000000; assign b = 64'h29B0000000000000;
    #10 assign a = 64'h130FFFFFFFFFFFFF; assign b = 64'h29BFFFFFFFFFFFFF;

    #10 $display("\n2**-718 * 2**-357:");
    #10 assign a = 64'h1310000000000000; assign b = 64'h29A0000000000000;
    #10 assign a = 64'h131FFFFFFFFFFFFF; assign b = 64'h29AFFFFFFFFFFFFF;

    #10 $display("\n2**-717 * 2**-358:");
    #10 assign a = 64'h1320000000000000; assign b = 64'h2990000000000000;
    #10 assign a = 64'h132FFFFFFFFFFFFF; assign b = 64'h299FFFFFFFFFFFFF;

    #10 $display("\n2**-716 * 2**-359:");
    #10 assign a = 64'h1330000000000000; assign b = 64'h2980000000000000;
    #10 assign a = 64'h133FFFFFFFFFFFFF; assign b = 64'h298FFFFFFFFFFFFF;

    #10 $display("\n2**-715 * 2**-360:");
    #10 assign a = 64'h1340000000000000; assign b = 64'h2970000000000000;
    #10 assign a = 64'h134FFFFFFFFFFFFF; assign b = 64'h297FFFFFFFFFFFFF;

    #10 $display("\n2**-714 * 2**-361:");
    #10 assign a = 64'h1350000000000000; assign b = 64'h2960000000000000;
    #10 assign a = 64'h135FFFFFFFFFFFFF; assign b = 64'h296FFFFFFFFFFFFF;

    #10 $display("\n2**-713 * 2**-362:");
    #10 assign a = 64'h1360000000000000; assign b = 64'h2950000000000000;
    #10 assign a = 64'h136FFFFFFFFFFFFF; assign b = 64'h295FFFFFFFFFFFFF;

    #10 $display("\n2**-712 * 2**-363:");
    #10 assign a = 64'h1370000000000000; assign b = 64'h2940000000000000;
    #10 assign a = 64'h137FFFFFFFFFFFFF; assign b = 64'h294FFFFFFFFFFFFF;

    #10 $display("\n2**-711 * 2**-364:");
    #10 assign a = 64'h1380000000000000; assign b = 64'h2930000000000000;
    #10 assign a = 64'h138FFFFFFFFFFFFF; assign b = 64'h293FFFFFFFFFFFFF;

    #10 $display("\n2**-710 * 2**-365:");
    #10 assign a = 64'h1390000000000000; assign b = 64'h2920000000000000;
    #10 assign a = 64'h139FFFFFFFFFFFFF; assign b = 64'h292FFFFFFFFFFFFF;

    #10 $display("\n2**-709 * 2**-366:");
    #10 assign a = 64'h13A0000000000000; assign b = 64'h2910000000000000;
    #10 assign a = 64'h13AFFFFFFFFFFFFF; assign b = 64'h291FFFFFFFFFFFFF;

    #10 $display("\n2**-708 * 2**-367:");
    #10 assign a = 64'h13B0000000000000; assign b = 64'h2900000000000000;
    #10 assign a = 64'h13BFFFFFFFFFFFFF; assign b = 64'h290FFFFFFFFFFFFF;

    #10 $display("\n2**-707 * 2**-368:");
    #10 assign a = 64'h13C0000000000000; assign b = 64'h28F0000000000000;
    #10 assign a = 64'h13CFFFFFFFFFFFFF; assign b = 64'h28FFFFFFFFFFFFFF;

    #10 $display("\n2**-706 * 2**-369:");
    #10 assign a = 64'h13D0000000000000; assign b = 64'h28E0000000000000;
    #10 assign a = 64'h13DFFFFFFFFFFFFF; assign b = 64'h28EFFFFFFFFFFFFF;

    #10 $display("\n2**-705 * 2**-370:");
    #10 assign a = 64'h13E0000000000000; assign b = 64'h28D0000000000000;
    #10 assign a = 64'h13EFFFFFFFFFFFFF; assign b = 64'h28DFFFFFFFFFFFFF;

    #10 $display("\n2**-704 * 2**-371:");
    #10 assign a = 64'h13F0000000000000; assign b = 64'h28C0000000000000;
    #10 assign a = 64'h13FFFFFFFFFFFFFF; assign b = 64'h28CFFFFFFFFFFFFF;

    #10 $display("\n2**-703 * 2**-372:");
    #10 assign a = 64'h1400000000000000; assign b = 64'h28B0000000000000;
    #10 assign a = 64'h140FFFFFFFFFFFFF; assign b = 64'h28BFFFFFFFFFFFFF;

    #10 $display("\n2**-702 * 2**-373:");
    #10 assign a = 64'h1410000000000000; assign b = 64'h28A0000000000000;
    #10 assign a = 64'h141FFFFFFFFFFFFF; assign b = 64'h28AFFFFFFFFFFFFF;

    #10 $display("\n2**-701 * 2**-374:");
    #10 assign a = 64'h1420000000000000; assign b = 64'h2890000000000000;
    #10 assign a = 64'h142FFFFFFFFFFFFF; assign b = 64'h289FFFFFFFFFFFFF;

    #10 $display("\n2**-700 * 2**-375:");
    #10 assign a = 64'h1430000000000000; assign b = 64'h2880000000000000;
    #10 assign a = 64'h143FFFFFFFFFFFFF; assign b = 64'h288FFFFFFFFFFFFF;

    #10 $display("\n2**-699 * 2**-376:");
    #10 assign a = 64'h1440000000000000; assign b = 64'h2870000000000000;
    #10 assign a = 64'h144FFFFFFFFFFFFF; assign b = 64'h287FFFFFFFFFFFFF;

    #10 $display("\n2**-698 * 2**-377:");
    #10 assign a = 64'h1450000000000000; assign b = 64'h2860000000000000;
    #10 assign a = 64'h145FFFFFFFFFFFFF; assign b = 64'h286FFFFFFFFFFFFF;

    #10 $display("\n2**-697 * 2**-378:");
    #10 assign a = 64'h1460000000000000; assign b = 64'h2850000000000000;
    #10 assign a = 64'h146FFFFFFFFFFFFF; assign b = 64'h285FFFFFFFFFFFFF;

    #10 $display("\n2**-696 * 2**-379:");
    #10 assign a = 64'h1470000000000000; assign b = 64'h2840000000000000;
    #10 assign a = 64'h147FFFFFFFFFFFFF; assign b = 64'h284FFFFFFFFFFFFF;

    #10 $display("\n2**-695 * 2**-380:");
    #10 assign a = 64'h1480000000000000; assign b = 64'h2830000000000000;
    #10 assign a = 64'h148FFFFFFFFFFFFF; assign b = 64'h283FFFFFFFFFFFFF;

    #10 $display("\n2**-694 * 2**-381:");
    #10 assign a = 64'h1490000000000000; assign b = 64'h2820000000000000;
    #10 assign a = 64'h149FFFFFFFFFFFFF; assign b = 64'h282FFFFFFFFFFFFF;

    #10 $display("\n2**-693 * 2**-382:");
    #10 assign a = 64'h14A0000000000000; assign b = 64'h2810000000000000;
    #10 assign a = 64'h14AFFFFFFFFFFFFF; assign b = 64'h281FFFFFFFFFFFFF;

    #10 $display("\n2**-692 * 2**-383:");
    #10 assign a = 64'h14B0000000000000; assign b = 64'h2800000000000000;
    #10 assign a = 64'h14BFFFFFFFFFFFFF; assign b = 64'h280FFFFFFFFFFFFF;

    #10 $display("\n2**-691 * 2**-384:");
    #10 assign a = 64'h14C0000000000000; assign b = 64'h27F0000000000000;
    #10 assign a = 64'h14CFFFFFFFFFFFFF; assign b = 64'h27FFFFFFFFFFFFFF;

    #10 $display("\n2**-690 * 2**-385:");
    #10 assign a = 64'h14D0000000000000; assign b = 64'h27E0000000000000;
    #10 assign a = 64'h14DFFFFFFFFFFFFF; assign b = 64'h27EFFFFFFFFFFFFF;

    #10 $display("\n2**-689 * 2**-386:");
    #10 assign a = 64'h14E0000000000000; assign b = 64'h27D0000000000000;
    #10 assign a = 64'h14EFFFFFFFFFFFFF; assign b = 64'h27DFFFFFFFFFFFFF;

    #10 $display("\n2**-688 * 2**-387:");
    #10 assign a = 64'h14F0000000000000; assign b = 64'h27C0000000000000;
    #10 assign a = 64'h14FFFFFFFFFFFFFF; assign b = 64'h27CFFFFFFFFFFFFF;

    #10 $display("\n2**-687 * 2**-388:");
    #10 assign a = 64'h1500000000000000; assign b = 64'h27B0000000000000;
    #10 assign a = 64'h150FFFFFFFFFFFFF; assign b = 64'h27BFFFFFFFFFFFFF;

    #10 $display("\n2**-686 * 2**-389:");
    #10 assign a = 64'h1510000000000000; assign b = 64'h27A0000000000000;
    #10 assign a = 64'h151FFFFFFFFFFFFF; assign b = 64'h27AFFFFFFFFFFFFF;

    #10 $display("\n2**-685 * 2**-390:");
    #10 assign a = 64'h1520000000000000; assign b = 64'h2790000000000000;
    #10 assign a = 64'h152FFFFFFFFFFFFF; assign b = 64'h279FFFFFFFFFFFFF;

    #10 $display("\n2**-684 * 2**-391:");
    #10 assign a = 64'h1530000000000000; assign b = 64'h2780000000000000;
    #10 assign a = 64'h153FFFFFFFFFFFFF; assign b = 64'h278FFFFFFFFFFFFF;

    #10 $display("\n2**-683 * 2**-392:");
    #10 assign a = 64'h1540000000000000; assign b = 64'h2770000000000000;
    #10 assign a = 64'h154FFFFFFFFFFFFF; assign b = 64'h277FFFFFFFFFFFFF;

    #10 $display("\n2**-682 * 2**-393:");
    #10 assign a = 64'h1550000000000000; assign b = 64'h2760000000000000;
    #10 assign a = 64'h155FFFFFFFFFFFFF; assign b = 64'h276FFFFFFFFFFFFF;

    #10 $display("\n2**-681 * 2**-394:");
    #10 assign a = 64'h1560000000000000; assign b = 64'h2750000000000000;
    #10 assign a = 64'h156FFFFFFFFFFFFF; assign b = 64'h275FFFFFFFFFFFFF;

    #10 $display("\n2**-680 * 2**-395:");
    #10 assign a = 64'h1570000000000000; assign b = 64'h2740000000000000;
    #10 assign a = 64'h157FFFFFFFFFFFFF; assign b = 64'h274FFFFFFFFFFFFF;

    #10 $display("\n2**-679 * 2**-396:");
    #10 assign a = 64'h1580000000000000; assign b = 64'h2730000000000000;
    #10 assign a = 64'h158FFFFFFFFFFFFF; assign b = 64'h273FFFFFFFFFFFFF;

    #10 $display("\n2**-678 * 2**-397:");
    #10 assign a = 64'h1590000000000000; assign b = 64'h2720000000000000;
    #10 assign a = 64'h159FFFFFFFFFFFFF; assign b = 64'h272FFFFFFFFFFFFF;

    #10 $display("\n2**-677 * 2**-398:");
    #10 assign a = 64'h15A0000000000000; assign b = 64'h2710000000000000;
    #10 assign a = 64'h15AFFFFFFFFFFFFF; assign b = 64'h271FFFFFFFFFFFFF;

    #10 $display("\n2**-676 * 2**-399:");
    #10 assign a = 64'h15B0000000000000; assign b = 64'h2700000000000000;
    #10 assign a = 64'h15BFFFFFFFFFFFFF; assign b = 64'h270FFFFFFFFFFFFF;

    #10 $display("\n2**-675 * 2**-400:");
    #10 assign a = 64'h15C0000000000000; assign b = 64'h26F0000000000000;
    #10 assign a = 64'h15CFFFFFFFFFFFFF; assign b = 64'h26FFFFFFFFFFFFFF;

    #10 $display("\n2**-674 * 2**-401:");
    #10 assign a = 64'h15D0000000000000; assign b = 64'h26E0000000000000;
    #10 assign a = 64'h15DFFFFFFFFFFFFF; assign b = 64'h26EFFFFFFFFFFFFF;

    #10 $display("\n2**-673 * 2**-402:");
    #10 assign a = 64'h15E0000000000000; assign b = 64'h26D0000000000000;
    #10 assign a = 64'h15EFFFFFFFFFFFFF; assign b = 64'h26DFFFFFFFFFFFFF;

    #10 $display("\n2**-672 * 2**-403:");
    #10 assign a = 64'h15F0000000000000; assign b = 64'h26C0000000000000;
    #10 assign a = 64'h15FFFFFFFFFFFFFF; assign b = 64'h26CFFFFFFFFFFFFF;

    #10 $display("\n2**-671 * 2**-404:");
    #10 assign a = 64'h1600000000000000; assign b = 64'h26B0000000000000;
    #10 assign a = 64'h160FFFFFFFFFFFFF; assign b = 64'h26BFFFFFFFFFFFFF;

    #10 $display("\n2**-670 * 2**-405:");
    #10 assign a = 64'h1610000000000000; assign b = 64'h26A0000000000000;
    #10 assign a = 64'h161FFFFFFFFFFFFF; assign b = 64'h26AFFFFFFFFFFFFF;

    #10 $display("\n2**-669 * 2**-406:");
    #10 assign a = 64'h1620000000000000; assign b = 64'h2690000000000000;
    #10 assign a = 64'h162FFFFFFFFFFFFF; assign b = 64'h269FFFFFFFFFFFFF;

    #10 $display("\n2**-668 * 2**-407:");
    #10 assign a = 64'h1630000000000000; assign b = 64'h2680000000000000;
    #10 assign a = 64'h163FFFFFFFFFFFFF; assign b = 64'h268FFFFFFFFFFFFF;

    #10 $display("\n2**-667 * 2**-408:");
    #10 assign a = 64'h1640000000000000; assign b = 64'h2670000000000000;
    #10 assign a = 64'h164FFFFFFFFFFFFF; assign b = 64'h267FFFFFFFFFFFFF;

    #10 $display("\n2**-666 * 2**-409:");
    #10 assign a = 64'h1650000000000000; assign b = 64'h2660000000000000;
    #10 assign a = 64'h165FFFFFFFFFFFFF; assign b = 64'h266FFFFFFFFFFFFF;

    #10 $display("\n2**-665 * 2**-410:");
    #10 assign a = 64'h1660000000000000; assign b = 64'h2650000000000000;
    #10 assign a = 64'h166FFFFFFFFFFFFF; assign b = 64'h265FFFFFFFFFFFFF;

    #10 $display("\n2**-664 * 2**-411:");
    #10 assign a = 64'h1670000000000000; assign b = 64'h2640000000000000;
    #10 assign a = 64'h167FFFFFFFFFFFFF; assign b = 64'h264FFFFFFFFFFFFF;

    #10 $display("\n2**-663 * 2**-412:");
    #10 assign a = 64'h1680000000000000; assign b = 64'h2630000000000000;
    #10 assign a = 64'h168FFFFFFFFFFFFF; assign b = 64'h263FFFFFFFFFFFFF;

    #10 $display("\n2**-662 * 2**-413:");
    #10 assign a = 64'h1690000000000000; assign b = 64'h2620000000000000;
    #10 assign a = 64'h169FFFFFFFFFFFFF; assign b = 64'h262FFFFFFFFFFFFF;

    #10 $display("\n2**-661 * 2**-414:");
    #10 assign a = 64'h16A0000000000000; assign b = 64'h2610000000000000;
    #10 assign a = 64'h16AFFFFFFFFFFFFF; assign b = 64'h261FFFFFFFFFFFFF;

    #10 $display("\n2**-660 * 2**-415:");
    #10 assign a = 64'h16B0000000000000; assign b = 64'h2600000000000000;
    #10 assign a = 64'h16BFFFFFFFFFFFFF; assign b = 64'h260FFFFFFFFFFFFF;

    #10 $display("\n2**-659 * 2**-416:");
    #10 assign a = 64'h16C0000000000000; assign b = 64'h25F0000000000000;
    #10 assign a = 64'h16CFFFFFFFFFFFFF; assign b = 64'h25FFFFFFFFFFFFFF;

    #10 $display("\n2**-658 * 2**-417:");
    #10 assign a = 64'h16D0000000000000; assign b = 64'h25E0000000000000;
    #10 assign a = 64'h16DFFFFFFFFFFFFF; assign b = 64'h25EFFFFFFFFFFFFF;

    #10 $display("\n2**-657 * 2**-418:");
    #10 assign a = 64'h16E0000000000000; assign b = 64'h25D0000000000000;
    #10 assign a = 64'h16EFFFFFFFFFFFFF; assign b = 64'h25DFFFFFFFFFFFFF;

    #10 $display("\n2**-656 * 2**-419:");
    #10 assign a = 64'h16F0000000000000; assign b = 64'h25C0000000000000;
    #10 assign a = 64'h16FFFFFFFFFFFFFF; assign b = 64'h25CFFFFFFFFFFFFF;

    #10 $display("\n2**-655 * 2**-420:");
    #10 assign a = 64'h1700000000000000; assign b = 64'h25B0000000000000;
    #10 assign a = 64'h170FFFFFFFFFFFFF; assign b = 64'h25BFFFFFFFFFFFFF;

    #10 $display("\n2**-654 * 2**-421:");
    #10 assign a = 64'h1710000000000000; assign b = 64'h25A0000000000000;
    #10 assign a = 64'h171FFFFFFFFFFFFF; assign b = 64'h25AFFFFFFFFFFFFF;

    #10 $display("\n2**-653 * 2**-422:");
    #10 assign a = 64'h1720000000000000; assign b = 64'h2590000000000000;
    #10 assign a = 64'h172FFFFFFFFFFFFF; assign b = 64'h259FFFFFFFFFFFFF;

    #10 $display("\n2**-652 * 2**-423:");
    #10 assign a = 64'h1730000000000000; assign b = 64'h2580000000000000;
    #10 assign a = 64'h173FFFFFFFFFFFFF; assign b = 64'h258FFFFFFFFFFFFF;

    #10 $display("\n2**-651 * 2**-424:");
    #10 assign a = 64'h1740000000000000; assign b = 64'h2570000000000000;
    #10 assign a = 64'h174FFFFFFFFFFFFF; assign b = 64'h257FFFFFFFFFFFFF;

    #10 $display("\n2**-650 * 2**-425:");
    #10 assign a = 64'h1750000000000000; assign b = 64'h2560000000000000;
    #10 assign a = 64'h175FFFFFFFFFFFFF; assign b = 64'h256FFFFFFFFFFFFF;

    #10 $display("\n2**-649 * 2**-426:");
    #10 assign a = 64'h1760000000000000; assign b = 64'h2550000000000000;
    #10 assign a = 64'h176FFFFFFFFFFFFF; assign b = 64'h255FFFFFFFFFFFFF;

    #10 $display("\n2**-648 * 2**-427:");
    #10 assign a = 64'h1770000000000000; assign b = 64'h2540000000000000;
    #10 assign a = 64'h177FFFFFFFFFFFFF; assign b = 64'h254FFFFFFFFFFFFF;

    #10 $display("\n2**-647 * 2**-428:");
    #10 assign a = 64'h1780000000000000; assign b = 64'h2530000000000000;
    #10 assign a = 64'h178FFFFFFFFFFFFF; assign b = 64'h253FFFFFFFFFFFFF;

    #10 $display("\n2**-646 * 2**-429:");
    #10 assign a = 64'h1790000000000000; assign b = 64'h2520000000000000;
    #10 assign a = 64'h179FFFFFFFFFFFFF; assign b = 64'h252FFFFFFFFFFFFF;

    #10 $display("\n2**-645 * 2**-430:");
    #10 assign a = 64'h17A0000000000000; assign b = 64'h2510000000000000;
    #10 assign a = 64'h17AFFFFFFFFFFFFF; assign b = 64'h251FFFFFFFFFFFFF;

    #10 $display("\n2**-644 * 2**-431:");
    #10 assign a = 64'h17B0000000000000; assign b = 64'h2500000000000000;
    #10 assign a = 64'h17BFFFFFFFFFFFFF; assign b = 64'h250FFFFFFFFFFFFF;

    #10 $display("\n2**-643 * 2**-432:");
    #10 assign a = 64'h17C0000000000000; assign b = 64'h24F0000000000000;
    #10 assign a = 64'h17CFFFFFFFFFFFFF; assign b = 64'h24FFFFFFFFFFFFFF;

    #10 $display("\n2**-642 * 2**-433:");
    #10 assign a = 64'h17D0000000000000; assign b = 64'h24E0000000000000;
    #10 assign a = 64'h17DFFFFFFFFFFFFF; assign b = 64'h24EFFFFFFFFFFFFF;

    #10 $display("\n2**-641 * 2**-434:");
    #10 assign a = 64'h17E0000000000000; assign b = 64'h24D0000000000000;
    #10 assign a = 64'h17EFFFFFFFFFFFFF; assign b = 64'h24DFFFFFFFFFFFFF;

    #10 $display("\n2**-640 * 2**-435:");
    #10 assign a = 64'h17F0000000000000; assign b = 64'h24C0000000000000;
    #10 assign a = 64'h17FFFFFFFFFFFFFF; assign b = 64'h24CFFFFFFFFFFFFF;

    #10 $display("\n2**-639 * 2**-436:");
    #10 assign a = 64'h1800000000000000; assign b = 64'h24B0000000000000;
    #10 assign a = 64'h180FFFFFFFFFFFFF; assign b = 64'h24BFFFFFFFFFFFFF;

    #10 $display("\n2**-638 * 2**-437:");
    #10 assign a = 64'h1810000000000000; assign b = 64'h24A0000000000000;
    #10 assign a = 64'h181FFFFFFFFFFFFF; assign b = 64'h24AFFFFFFFFFFFFF;

    #10 $display("\n2**-637 * 2**-438:");
    #10 assign a = 64'h1820000000000000; assign b = 64'h2490000000000000;
    #10 assign a = 64'h182FFFFFFFFFFFFF; assign b = 64'h249FFFFFFFFFFFFF;

    #10 $display("\n2**-636 * 2**-439:");
    #10 assign a = 64'h1830000000000000; assign b = 64'h2480000000000000;
    #10 assign a = 64'h183FFFFFFFFFFFFF; assign b = 64'h248FFFFFFFFFFFFF;

    #10 $display("\n2**-635 * 2**-440:");
    #10 assign a = 64'h1840000000000000; assign b = 64'h2470000000000000;
    #10 assign a = 64'h184FFFFFFFFFFFFF; assign b = 64'h247FFFFFFFFFFFFF;

    #10 $display("\n2**-634 * 2**-441:");
    #10 assign a = 64'h1850000000000000; assign b = 64'h2460000000000000;
    #10 assign a = 64'h185FFFFFFFFFFFFF; assign b = 64'h246FFFFFFFFFFFFF;

    #10 $display("\n2**-633 * 2**-442:");
    #10 assign a = 64'h1860000000000000; assign b = 64'h2450000000000000;
    #10 assign a = 64'h186FFFFFFFFFFFFF; assign b = 64'h245FFFFFFFFFFFFF;

    #10 $display("\n2**-632 * 2**-443:");
    #10 assign a = 64'h1870000000000000; assign b = 64'h2440000000000000;
    #10 assign a = 64'h187FFFFFFFFFFFFF; assign b = 64'h244FFFFFFFFFFFFF;

    #10 $display("\n2**-631 * 2**-444:");
    #10 assign a = 64'h1880000000000000; assign b = 64'h2430000000000000;
    #10 assign a = 64'h188FFFFFFFFFFFFF; assign b = 64'h243FFFFFFFFFFFFF;

    #10 $display("\n2**-630 * 2**-445:");
    #10 assign a = 64'h1890000000000000; assign b = 64'h2420000000000000;
    #10 assign a = 64'h189FFFFFFFFFFFFF; assign b = 64'h242FFFFFFFFFFFFF;

    #10 $display("\n2**-629 * 2**-446:");
    #10 assign a = 64'h18A0000000000000; assign b = 64'h2410000000000000;
    #10 assign a = 64'h18AFFFFFFFFFFFFF; assign b = 64'h241FFFFFFFFFFFFF;

    #10 $display("\n2**-628 * 2**-447:");
    #10 assign a = 64'h18B0000000000000; assign b = 64'h2400000000000000;
    #10 assign a = 64'h18BFFFFFFFFFFFFF; assign b = 64'h240FFFFFFFFFFFFF;

    #10 $display("\n2**-627 * 2**-448:");
    #10 assign a = 64'h18C0000000000000; assign b = 64'h23F0000000000000;
    #10 assign a = 64'h18CFFFFFFFFFFFFF; assign b = 64'h23FFFFFFFFFFFFFF;

    #10 $display("\n2**-626 * 2**-449:");
    #10 assign a = 64'h18D0000000000000; assign b = 64'h23E0000000000000;
    #10 assign a = 64'h18DFFFFFFFFFFFFF; assign b = 64'h23EFFFFFFFFFFFFF;

    #10 $display("\n2**-625 * 2**-450:");
    #10 assign a = 64'h18E0000000000000; assign b = 64'h23D0000000000000;
    #10 assign a = 64'h18EFFFFFFFFFFFFF; assign b = 64'h23DFFFFFFFFFFFFF;

    #10 $display("\n2**-624 * 2**-451:");
    #10 assign a = 64'h18F0000000000000; assign b = 64'h23C0000000000000;
    #10 assign a = 64'h18FFFFFFFFFFFFFF; assign b = 64'h23CFFFFFFFFFFFFF;

    #10 $display("\n2**-623 * 2**-452:");
    #10 assign a = 64'h1900000000000000; assign b = 64'h23B0000000000000;
    #10 assign a = 64'h190FFFFFFFFFFFFF; assign b = 64'h23BFFFFFFFFFFFFF;

    #10 $display("\n2**-622 * 2**-453:");
    #10 assign a = 64'h1910000000000000; assign b = 64'h23A0000000000000;
    #10 assign a = 64'h191FFFFFFFFFFFFF; assign b = 64'h23AFFFFFFFFFFFFF;

    #10 $display("\n2**-621 * 2**-454:");
    #10 assign a = 64'h1920000000000000; assign b = 64'h2390000000000000;
    #10 assign a = 64'h192FFFFFFFFFFFFF; assign b = 64'h239FFFFFFFFFFFFF;

    #10 $display("\n2**-620 * 2**-455:");
    #10 assign a = 64'h1930000000000000; assign b = 64'h2380000000000000;
    #10 assign a = 64'h193FFFFFFFFFFFFF; assign b = 64'h238FFFFFFFFFFFFF;

    #10 $display("\n2**-619 * 2**-456:");
    #10 assign a = 64'h1940000000000000; assign b = 64'h2370000000000000;
    #10 assign a = 64'h194FFFFFFFFFFFFF; assign b = 64'h237FFFFFFFFFFFFF;

    #10 $display("\n2**-618 * 2**-457:");
    #10 assign a = 64'h1950000000000000; assign b = 64'h2360000000000000;
    #10 assign a = 64'h195FFFFFFFFFFFFF; assign b = 64'h236FFFFFFFFFFFFF;

    #10 $display("\n2**-617 * 2**-458:");
    #10 assign a = 64'h1960000000000000; assign b = 64'h2350000000000000;
    #10 assign a = 64'h196FFFFFFFFFFFFF; assign b = 64'h235FFFFFFFFFFFFF;

    #10 $display("\n2**-616 * 2**-459:");
    #10 assign a = 64'h1970000000000000; assign b = 64'h2340000000000000;
    #10 assign a = 64'h197FFFFFFFFFFFFF; assign b = 64'h234FFFFFFFFFFFFF;

    #10 $display("\n2**-615 * 2**-460:");
    #10 assign a = 64'h1980000000000000; assign b = 64'h2330000000000000;
    #10 assign a = 64'h198FFFFFFFFFFFFF; assign b = 64'h233FFFFFFFFFFFFF;

    #10 $display("\n2**-614 * 2**-461:");
    #10 assign a = 64'h1990000000000000; assign b = 64'h2320000000000000;
    #10 assign a = 64'h199FFFFFFFFFFFFF; assign b = 64'h232FFFFFFFFFFFFF;

    #10 $display("\n2**-613 * 2**-462:");
    #10 assign a = 64'h19A0000000000000; assign b = 64'h2310000000000000;
    #10 assign a = 64'h19AFFFFFFFFFFFFF; assign b = 64'h231FFFFFFFFFFFFF;

    #10 $display("\n2**-612 * 2**-463:");
    #10 assign a = 64'h19B0000000000000; assign b = 64'h2300000000000000;
    #10 assign a = 64'h19BFFFFFFFFFFFFF; assign b = 64'h230FFFFFFFFFFFFF;

    #10 $display("\n2**-611 * 2**-464:");
    #10 assign a = 64'h19C0000000000000; assign b = 64'h22F0000000000000;
    #10 assign a = 64'h19CFFFFFFFFFFFFF; assign b = 64'h22FFFFFFFFFFFFFF;

    #10 $display("\n2**-610 * 2**-465:");
    #10 assign a = 64'h19D0000000000000; assign b = 64'h22E0000000000000;
    #10 assign a = 64'h19DFFFFFFFFFFFFF; assign b = 64'h22EFFFFFFFFFFFFF;

    #10 $display("\n2**-609 * 2**-466:");
    #10 assign a = 64'h19E0000000000000; assign b = 64'h22D0000000000000;
    #10 assign a = 64'h19EFFFFFFFFFFFFF; assign b = 64'h22DFFFFFFFFFFFFF;

    #10 $display("\n2**-608 * 2**-467:");
    #10 assign a = 64'h19F0000000000000; assign b = 64'h22C0000000000000;
    #10 assign a = 64'h19FFFFFFFFFFFFFF; assign b = 64'h22CFFFFFFFFFFFFF;

    #10 $display("\n2**-607 * 2**-468:");
    #10 assign a = 64'h1A00000000000000; assign b = 64'h22B0000000000000;
    #10 assign a = 64'h1A0FFFFFFFFFFFFF; assign b = 64'h22BFFFFFFFFFFFFF;

    #10 $display("\n2**-606 * 2**-469:");
    #10 assign a = 64'h1A10000000000000; assign b = 64'h22A0000000000000;
    #10 assign a = 64'h1A1FFFFFFFFFFFFF; assign b = 64'h22AFFFFFFFFFFFFF;

    #10 $display("\n2**-605 * 2**-470:");
    #10 assign a = 64'h1A20000000000000; assign b = 64'h2290000000000000;
    #10 assign a = 64'h1A2FFFFFFFFFFFFF; assign b = 64'h229FFFFFFFFFFFFF;

    #10 $display("\n2**-604 * 2**-471:");
    #10 assign a = 64'h1A30000000000000; assign b = 64'h2280000000000000;
    #10 assign a = 64'h1A3FFFFFFFFFFFFF; assign b = 64'h228FFFFFFFFFFFFF;

    #10 $display("\n2**-603 * 2**-472:");
    #10 assign a = 64'h1A40000000000000; assign b = 64'h2270000000000000;
    #10 assign a = 64'h1A4FFFFFFFFFFFFF; assign b = 64'h227FFFFFFFFFFFFF;

    #10 $display("\n2**-602 * 2**-473:");
    #10 assign a = 64'h1A50000000000000; assign b = 64'h2260000000000000;
    #10 assign a = 64'h1A5FFFFFFFFFFFFF; assign b = 64'h226FFFFFFFFFFFFF;

    #10 $display("\n2**-601 * 2**-474:");
    #10 assign a = 64'h1A60000000000000; assign b = 64'h2250000000000000;
    #10 assign a = 64'h1A6FFFFFFFFFFFFF; assign b = 64'h225FFFFFFFFFFFFF;

    #10 $display("\n2**-600 * 2**-475:");
    #10 assign a = 64'h1A70000000000000; assign b = 64'h2240000000000000;
    #10 assign a = 64'h1A7FFFFFFFFFFFFF; assign b = 64'h224FFFFFFFFFFFFF;

    #10 $display("\n2**-599 * 2**-476:");
    #10 assign a = 64'h1A80000000000000; assign b = 64'h2230000000000000;
    #10 assign a = 64'h1A8FFFFFFFFFFFFF; assign b = 64'h223FFFFFFFFFFFFF;

    #10 $display("\n2**-598 * 2**-477:");
    #10 assign a = 64'h1A90000000000000; assign b = 64'h2220000000000000;
    #10 assign a = 64'h1A9FFFFFFFFFFFFF; assign b = 64'h222FFFFFFFFFFFFF;

    #10 $display("\n2**-597 * 2**-478:");
    #10 assign a = 64'h1AA0000000000000; assign b = 64'h2210000000000000;
    #10 assign a = 64'h1AAFFFFFFFFFFFFF; assign b = 64'h221FFFFFFFFFFFFF;

    #10 $display("\n2**-596 * 2**-479:");
    #10 assign a = 64'h1AB0000000000000; assign b = 64'h2200000000000000;
    #10 assign a = 64'h1ABFFFFFFFFFFFFF; assign b = 64'h220FFFFFFFFFFFFF;

    #10 $display("\n2**-595 * 2**-480:");
    #10 assign a = 64'h1AC0000000000000; assign b = 64'h21F0000000000000;
    #10 assign a = 64'h1ACFFFFFFFFFFFFF; assign b = 64'h21FFFFFFFFFFFFFF;

    #10 $display("\n2**-594 * 2**-481:");
    #10 assign a = 64'h1AD0000000000000; assign b = 64'h21E0000000000000;
    #10 assign a = 64'h1ADFFFFFFFFFFFFF; assign b = 64'h21EFFFFFFFFFFFFF;

    #10 $display("\n2**-593 * 2**-482:");
    #10 assign a = 64'h1AE0000000000000; assign b = 64'h21D0000000000000;
    #10 assign a = 64'h1AEFFFFFFFFFFFFF; assign b = 64'h21DFFFFFFFFFFFFF;

    #10 $display("\n2**-592 * 2**-483:");
    #10 assign a = 64'h1AF0000000000000; assign b = 64'h21C0000000000000;
    #10 assign a = 64'h1AFFFFFFFFFFFFFF; assign b = 64'h21CFFFFFFFFFFFFF;

    #10 $display("\n2**-591 * 2**-484:");
    #10 assign a = 64'h1B00000000000000; assign b = 64'h21B0000000000000;
    #10 assign a = 64'h1B0FFFFFFFFFFFFF; assign b = 64'h21BFFFFFFFFFFFFF;

    #10 $display("\n2**-590 * 2**-485:");
    #10 assign a = 64'h1B10000000000000; assign b = 64'h21A0000000000000;
    #10 assign a = 64'h1B1FFFFFFFFFFFFF; assign b = 64'h21AFFFFFFFFFFFFF;

    #10 $display("\n2**-589 * 2**-486:");
    #10 assign a = 64'h1B20000000000000; assign b = 64'h2190000000000000;
    #10 assign a = 64'h1B2FFFFFFFFFFFFF; assign b = 64'h219FFFFFFFFFFFFF;

    #10 $display("\n2**-588 * 2**-487:");
    #10 assign a = 64'h1B30000000000000; assign b = 64'h2180000000000000;
    #10 assign a = 64'h1B3FFFFFFFFFFFFF; assign b = 64'h218FFFFFFFFFFFFF;

    #10 $display("\n2**-587 * 2**-488:");
    #10 assign a = 64'h1B40000000000000; assign b = 64'h2170000000000000;
    #10 assign a = 64'h1B4FFFFFFFFFFFFF; assign b = 64'h217FFFFFFFFFFFFF;

    #10 $display("\n2**-586 * 2**-489:");
    #10 assign a = 64'h1B50000000000000; assign b = 64'h2160000000000000;
    #10 assign a = 64'h1B5FFFFFFFFFFFFF; assign b = 64'h216FFFFFFFFFFFFF;

    #10 $display("\n2**-585 * 2**-490:");
    #10 assign a = 64'h1B60000000000000; assign b = 64'h2150000000000000;
    #10 assign a = 64'h1B6FFFFFFFFFFFFF; assign b = 64'h215FFFFFFFFFFFFF;

    #10 $display("\n2**-584 * 2**-491:");
    #10 assign a = 64'h1B70000000000000; assign b = 64'h2140000000000000;
    #10 assign a = 64'h1B7FFFFFFFFFFFFF; assign b = 64'h214FFFFFFFFFFFFF;

    #10 $display("\n2**-583 * 2**-492:");
    #10 assign a = 64'h1B80000000000000; assign b = 64'h2130000000000000;
    #10 assign a = 64'h1B8FFFFFFFFFFFFF; assign b = 64'h213FFFFFFFFFFFFF;

    #10 $display("\n2**-582 * 2**-493:");
    #10 assign a = 64'h1B90000000000000; assign b = 64'h2120000000000000;
    #10 assign a = 64'h1B9FFFFFFFFFFFFF; assign b = 64'h212FFFFFFFFFFFFF;

    #10 $display("\n2**-581 * 2**-494:");
    #10 assign a = 64'h1BA0000000000000; assign b = 64'h2110000000000000;
    #10 assign a = 64'h1BAFFFFFFFFFFFFF; assign b = 64'h211FFFFFFFFFFFFF;

    #10 $display("\n2**-580 * 2**-495:");
    #10 assign a = 64'h1BB0000000000000; assign b = 64'h2100000000000000;
    #10 assign a = 64'h1BBFFFFFFFFFFFFF; assign b = 64'h210FFFFFFFFFFFFF;

    #10 $display("\n2**-579 * 2**-496:");
    #10 assign a = 64'h1BC0000000000000; assign b = 64'h20F0000000000000;
    #10 assign a = 64'h1BCFFFFFFFFFFFFF; assign b = 64'h20FFFFFFFFFFFFFF;

    #10 $display("\n2**-578 * 2**-497:");
    #10 assign a = 64'h1BD0000000000000; assign b = 64'h20E0000000000000;
    #10 assign a = 64'h1BDFFFFFFFFFFFFF; assign b = 64'h20EFFFFFFFFFFFFF;

    #10 $display("\n2**-577 * 2**-498:");
    #10 assign a = 64'h1BE0000000000000; assign b = 64'h20D0000000000000;
    #10 assign a = 64'h1BEFFFFFFFFFFFFF; assign b = 64'h20DFFFFFFFFFFFFF;

    #10 $display("\n2**-576 * 2**-499:");
    #10 assign a = 64'h1BF0000000000000; assign b = 64'h20C0000000000000;
    #10 assign a = 64'h1BFFFFFFFFFFFFFF; assign b = 64'h20CFFFFFFFFFFFFF;

    #10 $display("\n2**-575 * 2**-500:");
    #10 assign a = 64'h1C00000000000000; assign b = 64'h20B0000000000000;
    #10 assign a = 64'h1C0FFFFFFFFFFFFF; assign b = 64'h20BFFFFFFFFFFFFF;

    #10 $display("\n2**-574 * 2**-501:");
    #10 assign a = 64'h1C10000000000000; assign b = 64'h20A0000000000000;
    #10 assign a = 64'h1C1FFFFFFFFFFFFF; assign b = 64'h20AFFFFFFFFFFFFF;

    #10 $display("\n2**-573 * 2**-502:");
    #10 assign a = 64'h1C20000000000000; assign b = 64'h2090000000000000;
    #10 assign a = 64'h1C2FFFFFFFFFFFFF; assign b = 64'h209FFFFFFFFFFFFF;

    #10 $display("\n2**-572 * 2**-503:");
    #10 assign a = 64'h1C30000000000000; assign b = 64'h2080000000000000;
    #10 assign a = 64'h1C3FFFFFFFFFFFFF; assign b = 64'h208FFFFFFFFFFFFF;

    #10 $display("\n2**-571 * 2**-504:");
    #10 assign a = 64'h1C40000000000000; assign b = 64'h2070000000000000;
    #10 assign a = 64'h1C4FFFFFFFFFFFFF; assign b = 64'h207FFFFFFFFFFFFF;

    #10 $display("\n2**-570 * 2**-505:");
    #10 assign a = 64'h1C50000000000000; assign b = 64'h2060000000000000;
    #10 assign a = 64'h1C5FFFFFFFFFFFFF; assign b = 64'h206FFFFFFFFFFFFF;

    #10 $display("\n2**-569 * 2**-506:");
    #10 assign a = 64'h1C60000000000000; assign b = 64'h2050000000000000;
    #10 assign a = 64'h1C6FFFFFFFFFFFFF; assign b = 64'h205FFFFFFFFFFFFF;

    #10 $display("\n2**-568 * 2**-507:");
    #10 assign a = 64'h1C70000000000000; assign b = 64'h2040000000000000;
    #10 assign a = 64'h1C7FFFFFFFFFFFFF; assign b = 64'h204FFFFFFFFFFFFF;

    #10 $display("\n2**-567 * 2**-508:");
    #10 assign a = 64'h1C80000000000000; assign b = 64'h2030000000000000;
    #10 assign a = 64'h1C8FFFFFFFFFFFFF; assign b = 64'h203FFFFFFFFFFFFF;

    #10 $display("\n2**-566 * 2**-509:");
    #10 assign a = 64'h1C90000000000000; assign b = 64'h2020000000000000;
    #10 assign a = 64'h1C9FFFFFFFFFFFFF; assign b = 64'h202FFFFFFFFFFFFF;

    #10 $display("\n2**-565 * 2**-510:");
    #10 assign a = 64'h1CA0000000000000; assign b = 64'h2010000000000000;
    #10 assign a = 64'h1CAFFFFFFFFFFFFF; assign b = 64'h201FFFFFFFFFFFFF;

    #10 $display("\n2**-564 * 2**-511:");
    #10 assign a = 64'h1CB0000000000000; assign b = 64'h2000000000000000;
    #10 assign a = 64'h1CBFFFFFFFFFFFFF; assign b = 64'h200FFFFFFFFFFFFF;

    #10 $display("\n2**-563 * 2**-512:");
    #10 assign a = 64'h1CC0000000000000; assign b = 64'h1FF0000000000000;
    #10 assign a = 64'h1CCFFFFFFFFFFFFF; assign b = 64'h1FFFFFFFFFFFFFFF;

    #10 $display("\n2**-562 * 2**-513:");
    #10 assign a = 64'h1CD0000000000000; assign b = 64'h1FE0000000000000;
    #10 assign a = 64'h1CDFFFFFFFFFFFFF; assign b = 64'h1FEFFFFFFFFFFFFF;

    #10 $display("\n2**-561 * 2**-514:");
    #10 assign a = 64'h1CE0000000000000; assign b = 64'h1FD0000000000000;
    #10 assign a = 64'h1CEFFFFFFFFFFFFF; assign b = 64'h1FDFFFFFFFFFFFFF;

    #10 $display("\n2**-560 * 2**-515:");
    #10 assign a = 64'h1CF0000000000000; assign b = 64'h1FC0000000000000;
    #10 assign a = 64'h1CFFFFFFFFFFFFFF; assign b = 64'h1FCFFFFFFFFFFFFF;

    #10 $display("\n2**-559 * 2**-516:");
    #10 assign a = 64'h1D00000000000000; assign b = 64'h1FB0000000000000;
    #10 assign a = 64'h1D0FFFFFFFFFFFFF; assign b = 64'h1FBFFFFFFFFFFFFF;

    #10 $display("\n2**-558 * 2**-517:");
    #10 assign a = 64'h1D10000000000000; assign b = 64'h1FA0000000000000;
    #10 assign a = 64'h1D1FFFFFFFFFFFFF; assign b = 64'h1FAFFFFFFFFFFFFF;

    #10 $display("\n2**-557 * 2**-518:");
    #10 assign a = 64'h1D20000000000000; assign b = 64'h1F90000000000000;
    #10 assign a = 64'h1D2FFFFFFFFFFFFF; assign b = 64'h1F9FFFFFFFFFFFFF;

    #10 $display("\n2**-556 * 2**-519:");
    #10 assign a = 64'h1D30000000000000; assign b = 64'h1F80000000000000;
    #10 assign a = 64'h1D3FFFFFFFFFFFFF; assign b = 64'h1F8FFFFFFFFFFFFF;

    #10 $display("\n2**-555 * 2**-520:");
    #10 assign a = 64'h1D40000000000000; assign b = 64'h1F70000000000000;
    #10 assign a = 64'h1D4FFFFFFFFFFFFF; assign b = 64'h1F7FFFFFFFFFFFFF;

    #10 $display("\n2**-554 * 2**-521:");
    #10 assign a = 64'h1D50000000000000; assign b = 64'h1F60000000000000;
    #10 assign a = 64'h1D5FFFFFFFFFFFFF; assign b = 64'h1F6FFFFFFFFFFFFF;

    #10 $display("\n2**-553 * 2**-522:");
    #10 assign a = 64'h1D60000000000000; assign b = 64'h1F50000000000000;
    #10 assign a = 64'h1D6FFFFFFFFFFFFF; assign b = 64'h1F5FFFFFFFFFFFFF;

    #10 $display("\n2**-552 * 2**-523:");
    #10 assign a = 64'h1D70000000000000; assign b = 64'h1F40000000000000;
    #10 assign a = 64'h1D7FFFFFFFFFFFFF; assign b = 64'h1F4FFFFFFFFFFFFF;

    #10 $display("\n2**-551 * 2**-524:");
    #10 assign a = 64'h1D80000000000000; assign b = 64'h1F30000000000000;
    #10 assign a = 64'h1D8FFFFFFFFFFFFF; assign b = 64'h1F3FFFFFFFFFFFFF;

    #10 $display("\n2**-550 * 2**-525:");
    #10 assign a = 64'h1D90000000000000; assign b = 64'h1F20000000000000;
    #10 assign a = 64'h1D9FFFFFFFFFFFFF; assign b = 64'h1F2FFFFFFFFFFFFF;

    #10 $display("\n2**-549 * 2**-526:");
    #10 assign a = 64'h1DA0000000000000; assign b = 64'h1F10000000000000;
    #10 assign a = 64'h1DAFFFFFFFFFFFFF; assign b = 64'h1F1FFFFFFFFFFFFF;

    #10 $display("\n2**-548 * 2**-527:");
    #10 assign a = 64'h1DB0000000000000; assign b = 64'h1F00000000000000;
    #10 assign a = 64'h1DBFFFFFFFFFFFFF; assign b = 64'h1F0FFFFFFFFFFFFF;

    #10 $display("\n2**-547 * 2**-528:");
    #10 assign a = 64'h1DC0000000000000; assign b = 64'h1EF0000000000000;
    #10 assign a = 64'h1DCFFFFFFFFFFFFF; assign b = 64'h1EFFFFFFFFFFFFFF;

    #10 $display("\n2**-546 * 2**-529:");
    #10 assign a = 64'h1DD0000000000000; assign b = 64'h1EE0000000000000;
    #10 assign a = 64'h1DDFFFFFFFFFFFFF; assign b = 64'h1EEFFFFFFFFFFFFF;

    #10 $display("\n2**-545 * 2**-530:");
    #10 assign a = 64'h1DE0000000000000; assign b = 64'h1ED0000000000000;
    #10 assign a = 64'h1DEFFFFFFFFFFFFF; assign b = 64'h1EDFFFFFFFFFFFFF;

    #10 $display("\n2**-544 * 2**-531:");
    #10 assign a = 64'h1DF0000000000000; assign b = 64'h1EC0000000000000;
    #10 assign a = 64'h1DFFFFFFFFFFFFFF; assign b = 64'h1ECFFFFFFFFFFFFF;

    #10 $display("\n2**-543 * 2**-532:");
    #10 assign a = 64'h1E00000000000000; assign b = 64'h1EB0000000000000;
    #10 assign a = 64'h1E0FFFFFFFFFFFFF; assign b = 64'h1EBFFFFFFFFFFFFF;

    #10 $display("\n2**-542 * 2**-533:");
    #10 assign a = 64'h1E10000000000000; assign b = 64'h1EA0000000000000;
    #10 assign a = 64'h1E1FFFFFFFFFFFFF; assign b = 64'h1EAFFFFFFFFFFFFF;

    #10 $display("\n2**-541 * 2**-534:");
    #10 assign a = 64'h1E20000000000000; assign b = 64'h1E90000000000000;
    #10 assign a = 64'h1E2FFFFFFFFFFFFF; assign b = 64'h1E9FFFFFFFFFFFFF;

    #10 $display("\n2**-540 * 2**-535:");
    #10 assign a = 64'h1E30000000000000; assign b = 64'h1E80000000000000;
    #10 assign a = 64'h1E3FFFFFFFFFFFFF; assign b = 64'h1E8FFFFFFFFFFFFF;

    #10 $display("\n2**-539 * 2**-536:");
    #10 assign a = 64'h1E40000000000000; assign b = 64'h1E70000000000000;
    #10 assign a = 64'h1E4FFFFFFFFFFFFF; assign b = 64'h1E7FFFFFFFFFFFFF;

    #10 $display("\n2**-538 * 2**-537:");
    #10 assign a = 64'h1E50000000000000; assign b = 64'h1E60000000000000;
    #10 assign a = 64'h1E5FFFFFFFFFFFFF; assign b = 64'h1E6FFFFFFFFFFFFF;

    #10 $display("\n2**-537 * 2**-538:");
    #10 assign a = 64'h1E60000000000000; assign b = 64'h1E50000000000000;
    #10 assign a = 64'h1E6FFFFFFFFFFFFF; assign b = 64'h1E5FFFFFFFFFFFFF;

    #10 $display("\n2**-536 * 2**-539:");
    #10 assign a = 64'h1E70000000000000; assign b = 64'h1E40000000000000;
    #10 assign a = 64'h1E7FFFFFFFFFFFFF; assign b = 64'h1E4FFFFFFFFFFFFF;

    #10 $display("\n2**-535 * 2**-540:");
    #10 assign a = 64'h1E80000000000000; assign b = 64'h1E30000000000000;
    #10 assign a = 64'h1E8FFFFFFFFFFFFF; assign b = 64'h1E3FFFFFFFFFFFFF;

    #10 $display("\n2**-534 * 2**-541:");
    #10 assign a = 64'h1E90000000000000; assign b = 64'h1E20000000000000;
    #10 assign a = 64'h1E9FFFFFFFFFFFFF; assign b = 64'h1E2FFFFFFFFFFFFF;

    #10 $display("\n2**-533 * 2**-542:");
    #10 assign a = 64'h1EA0000000000000; assign b = 64'h1E10000000000000;
    #10 assign a = 64'h1EAFFFFFFFFFFFFF; assign b = 64'h1E1FFFFFFFFFFFFF;

    #10 $display("\n2**-532 * 2**-543:");
    #10 assign a = 64'h1EB0000000000000; assign b = 64'h1E00000000000000;
    #10 assign a = 64'h1EBFFFFFFFFFFFFF; assign b = 64'h1E0FFFFFFFFFFFFF;

    #10 $display("\n2**-531 * 2**-544:");
    #10 assign a = 64'h1EC0000000000000; assign b = 64'h1DF0000000000000;
    #10 assign a = 64'h1ECFFFFFFFFFFFFF; assign b = 64'h1DFFFFFFFFFFFFFF;

    #10 $display("\n2**-530 * 2**-545:");
    #10 assign a = 64'h1ED0000000000000; assign b = 64'h1DE0000000000000;
    #10 assign a = 64'h1EDFFFFFFFFFFFFF; assign b = 64'h1DEFFFFFFFFFFFFF;

    #10 $display("\n2**-529 * 2**-546:");
    #10 assign a = 64'h1EE0000000000000; assign b = 64'h1DD0000000000000;
    #10 assign a = 64'h1EEFFFFFFFFFFFFF; assign b = 64'h1DDFFFFFFFFFFFFF;

    #10 $display("\n2**-528 * 2**-547:");
    #10 assign a = 64'h1EF0000000000000; assign b = 64'h1DC0000000000000;
    #10 assign a = 64'h1EFFFFFFFFFFFFFF; assign b = 64'h1DCFFFFFFFFFFFFF;

    #10 $display("\n2**-527 * 2**-548:");
    #10 assign a = 64'h1F00000000000000; assign b = 64'h1DB0000000000000;
    #10 assign a = 64'h1F0FFFFFFFFFFFFF; assign b = 64'h1DBFFFFFFFFFFFFF;

    #10 $display("\n2**-526 * 2**-549:");
    #10 assign a = 64'h1F10000000000000; assign b = 64'h1DA0000000000000;
    #10 assign a = 64'h1F1FFFFFFFFFFFFF; assign b = 64'h1DAFFFFFFFFFFFFF;

    #10 $display("\n2**-525 * 2**-550:");
    #10 assign a = 64'h1F20000000000000; assign b = 64'h1D90000000000000;
    #10 assign a = 64'h1F2FFFFFFFFFFFFF; assign b = 64'h1D9FFFFFFFFFFFFF;

    #10 $display("\n2**-524 * 2**-551:");
    #10 assign a = 64'h1F30000000000000; assign b = 64'h1D80000000000000;
    #10 assign a = 64'h1F3FFFFFFFFFFFFF; assign b = 64'h1D8FFFFFFFFFFFFF;

    #10 $display("\n2**-523 * 2**-552:");
    #10 assign a = 64'h1F40000000000000; assign b = 64'h1D70000000000000;
    #10 assign a = 64'h1F4FFFFFFFFFFFFF; assign b = 64'h1D7FFFFFFFFFFFFF;

    #10 $display("\n2**-522 * 2**-553:");
    #10 assign a = 64'h1F50000000000000; assign b = 64'h1D60000000000000;
    #10 assign a = 64'h1F5FFFFFFFFFFFFF; assign b = 64'h1D6FFFFFFFFFFFFF;

    #10 $display("\n2**-521 * 2**-554:");
    #10 assign a = 64'h1F60000000000000; assign b = 64'h1D50000000000000;
    #10 assign a = 64'h1F6FFFFFFFFFFFFF; assign b = 64'h1D5FFFFFFFFFFFFF;

    #10 $display("\n2**-520 * 2**-555:");
    #10 assign a = 64'h1F70000000000000; assign b = 64'h1D40000000000000;
    #10 assign a = 64'h1F7FFFFFFFFFFFFF; assign b = 64'h1D4FFFFFFFFFFFFF;

    #10 $display("\n2**-519 * 2**-556:");
    #10 assign a = 64'h1F80000000000000; assign b = 64'h1D30000000000000;
    #10 assign a = 64'h1F8FFFFFFFFFFFFF; assign b = 64'h1D3FFFFFFFFFFFFF;

    #10 $display("\n2**-518 * 2**-557:");
    #10 assign a = 64'h1F90000000000000; assign b = 64'h1D20000000000000;
    #10 assign a = 64'h1F9FFFFFFFFFFFFF; assign b = 64'h1D2FFFFFFFFFFFFF;

    #10 $display("\n2**-517 * 2**-558:");
    #10 assign a = 64'h1FA0000000000000; assign b = 64'h1D10000000000000;
    #10 assign a = 64'h1FAFFFFFFFFFFFFF; assign b = 64'h1D1FFFFFFFFFFFFF;

    #10 $display("\n2**-516 * 2**-559:");
    #10 assign a = 64'h1FB0000000000000; assign b = 64'h1D00000000000000;
    #10 assign a = 64'h1FBFFFFFFFFFFFFF; assign b = 64'h1D0FFFFFFFFFFFFF;

    #10 $display("\n2**-515 * 2**-560:");
    #10 assign a = 64'h1FC0000000000000; assign b = 64'h1CF0000000000000;
    #10 assign a = 64'h1FCFFFFFFFFFFFFF; assign b = 64'h1CFFFFFFFFFFFFFF;

    #10 $display("\n2**-514 * 2**-561:");
    #10 assign a = 64'h1FD0000000000000; assign b = 64'h1CE0000000000000;
    #10 assign a = 64'h1FDFFFFFFFFFFFFF; assign b = 64'h1CEFFFFFFFFFFFFF;

    #10 $display("\n2**-513 * 2**-562:");
    #10 assign a = 64'h1FE0000000000000; assign b = 64'h1CD0000000000000;
    #10 assign a = 64'h1FEFFFFFFFFFFFFF; assign b = 64'h1CDFFFFFFFFFFFFF;

    #10 $display("\n2**-512 * 2**-563:");
    #10 assign a = 64'h1FF0000000000000; assign b = 64'h1CC0000000000000;
    #10 assign a = 64'h1FFFFFFFFFFFFFFF; assign b = 64'h1CCFFFFFFFFFFFFF;

    #10 $display("\n2**-511 * 2**-564:");
    #10 assign a = 64'h2000000000000000; assign b = 64'h1CB0000000000000;
    #10 assign a = 64'h200FFFFFFFFFFFFF; assign b = 64'h1CBFFFFFFFFFFFFF;

    #10 $display("\n2**-510 * 2**-565:");
    #10 assign a = 64'h2010000000000000; assign b = 64'h1CA0000000000000;
    #10 assign a = 64'h201FFFFFFFFFFFFF; assign b = 64'h1CAFFFFFFFFFFFFF;

    #10 $display("\n2**-509 * 2**-566:");
    #10 assign a = 64'h2020000000000000; assign b = 64'h1C90000000000000;
    #10 assign a = 64'h202FFFFFFFFFFFFF; assign b = 64'h1C9FFFFFFFFFFFFF;

    #10 $display("\n2**-508 * 2**-567:");
    #10 assign a = 64'h2030000000000000; assign b = 64'h1C80000000000000;
    #10 assign a = 64'h203FFFFFFFFFFFFF; assign b = 64'h1C8FFFFFFFFFFFFF;

    #10 $display("\n2**-507 * 2**-568:");
    #10 assign a = 64'h2040000000000000; assign b = 64'h1C70000000000000;
    #10 assign a = 64'h204FFFFFFFFFFFFF; assign b = 64'h1C7FFFFFFFFFFFFF;

    #10 $display("\n2**-506 * 2**-569:");
    #10 assign a = 64'h2050000000000000; assign b = 64'h1C60000000000000;
    #10 assign a = 64'h205FFFFFFFFFFFFF; assign b = 64'h1C6FFFFFFFFFFFFF;

    #10 $display("\n2**-505 * 2**-570:");
    #10 assign a = 64'h2060000000000000; assign b = 64'h1C50000000000000;
    #10 assign a = 64'h206FFFFFFFFFFFFF; assign b = 64'h1C5FFFFFFFFFFFFF;

    #10 $display("\n2**-504 * 2**-571:");
    #10 assign a = 64'h2070000000000000; assign b = 64'h1C40000000000000;
    #10 assign a = 64'h207FFFFFFFFFFFFF; assign b = 64'h1C4FFFFFFFFFFFFF;

    #10 $display("\n2**-503 * 2**-572:");
    #10 assign a = 64'h2080000000000000; assign b = 64'h1C30000000000000;
    #10 assign a = 64'h208FFFFFFFFFFFFF; assign b = 64'h1C3FFFFFFFFFFFFF;

    #10 $display("\n2**-502 * 2**-573:");
    #10 assign a = 64'h2090000000000000; assign b = 64'h1C20000000000000;
    #10 assign a = 64'h209FFFFFFFFFFFFF; assign b = 64'h1C2FFFFFFFFFFFFF;

    #10 $display("\n2**-501 * 2**-574:");
    #10 assign a = 64'h20A0000000000000; assign b = 64'h1C10000000000000;
    #10 assign a = 64'h20AFFFFFFFFFFFFF; assign b = 64'h1C1FFFFFFFFFFFFF;

    #10 $display("\n2**-500 * 2**-575:");
    #10 assign a = 64'h20B0000000000000; assign b = 64'h1C00000000000000;
    #10 assign a = 64'h20BFFFFFFFFFFFFF; assign b = 64'h1C0FFFFFFFFFFFFF;

    #10 $display("\n2**-499 * 2**-576:");
    #10 assign a = 64'h20C0000000000000; assign b = 64'h1BF0000000000000;
    #10 assign a = 64'h20CFFFFFFFFFFFFF; assign b = 64'h1BFFFFFFFFFFFFFF;

    #10 $display("\n2**-498 * 2**-577:");
    #10 assign a = 64'h20D0000000000000; assign b = 64'h1BE0000000000000;
    #10 assign a = 64'h20DFFFFFFFFFFFFF; assign b = 64'h1BEFFFFFFFFFFFFF;

    #10 $display("\n2**-497 * 2**-578:");
    #10 assign a = 64'h20E0000000000000; assign b = 64'h1BD0000000000000;
    #10 assign a = 64'h20EFFFFFFFFFFFFF; assign b = 64'h1BDFFFFFFFFFFFFF;

    #10 $display("\n2**-496 * 2**-579:");
    #10 assign a = 64'h20F0000000000000; assign b = 64'h1BC0000000000000;
    #10 assign a = 64'h20FFFFFFFFFFFFFF; assign b = 64'h1BCFFFFFFFFFFFFF;

    #10 $display("\n2**-495 * 2**-580:");
    #10 assign a = 64'h2100000000000000; assign b = 64'h1BB0000000000000;
    #10 assign a = 64'h210FFFFFFFFFFFFF; assign b = 64'h1BBFFFFFFFFFFFFF;

    #10 $display("\n2**-494 * 2**-581:");
    #10 assign a = 64'h2110000000000000; assign b = 64'h1BA0000000000000;
    #10 assign a = 64'h211FFFFFFFFFFFFF; assign b = 64'h1BAFFFFFFFFFFFFF;

    #10 $display("\n2**-493 * 2**-582:");
    #10 assign a = 64'h2120000000000000; assign b = 64'h1B90000000000000;
    #10 assign a = 64'h212FFFFFFFFFFFFF; assign b = 64'h1B9FFFFFFFFFFFFF;

    #10 $display("\n2**-492 * 2**-583:");
    #10 assign a = 64'h2130000000000000; assign b = 64'h1B80000000000000;
    #10 assign a = 64'h213FFFFFFFFFFFFF; assign b = 64'h1B8FFFFFFFFFFFFF;

    #10 $display("\n2**-491 * 2**-584:");
    #10 assign a = 64'h2140000000000000; assign b = 64'h1B70000000000000;
    #10 assign a = 64'h214FFFFFFFFFFFFF; assign b = 64'h1B7FFFFFFFFFFFFF;

    #10 $display("\n2**-490 * 2**-585:");
    #10 assign a = 64'h2150000000000000; assign b = 64'h1B60000000000000;
    #10 assign a = 64'h215FFFFFFFFFFFFF; assign b = 64'h1B6FFFFFFFFFFFFF;

    #10 $display("\n2**-489 * 2**-586:");
    #10 assign a = 64'h2160000000000000; assign b = 64'h1B50000000000000;
    #10 assign a = 64'h216FFFFFFFFFFFFF; assign b = 64'h1B5FFFFFFFFFFFFF;

    #10 $display("\n2**-488 * 2**-587:");
    #10 assign a = 64'h2170000000000000; assign b = 64'h1B40000000000000;
    #10 assign a = 64'h217FFFFFFFFFFFFF; assign b = 64'h1B4FFFFFFFFFFFFF;

    #10 $display("\n2**-487 * 2**-588:");
    #10 assign a = 64'h2180000000000000; assign b = 64'h1B30000000000000;
    #10 assign a = 64'h218FFFFFFFFFFFFF; assign b = 64'h1B3FFFFFFFFFFFFF;

    #10 $display("\n2**-486 * 2**-589:");
    #10 assign a = 64'h2190000000000000; assign b = 64'h1B20000000000000;
    #10 assign a = 64'h219FFFFFFFFFFFFF; assign b = 64'h1B2FFFFFFFFFFFFF;

    #10 $display("\n2**-485 * 2**-590:");
    #10 assign a = 64'h21A0000000000000; assign b = 64'h1B10000000000000;
    #10 assign a = 64'h21AFFFFFFFFFFFFF; assign b = 64'h1B1FFFFFFFFFFFFF;

    #10 $display("\n2**-484 * 2**-591:");
    #10 assign a = 64'h21B0000000000000; assign b = 64'h1B00000000000000;
    #10 assign a = 64'h21BFFFFFFFFFFFFF; assign b = 64'h1B0FFFFFFFFFFFFF;

    #10 $display("\n2**-483 * 2**-592:");
    #10 assign a = 64'h21C0000000000000; assign b = 64'h1AF0000000000000;
    #10 assign a = 64'h21CFFFFFFFFFFFFF; assign b = 64'h1AFFFFFFFFFFFFFF;

    #10 $display("\n2**-482 * 2**-593:");
    #10 assign a = 64'h21D0000000000000; assign b = 64'h1AE0000000000000;
    #10 assign a = 64'h21DFFFFFFFFFFFFF; assign b = 64'h1AEFFFFFFFFFFFFF;

    #10 $display("\n2**-481 * 2**-594:");
    #10 assign a = 64'h21E0000000000000; assign b = 64'h1AD0000000000000;
    #10 assign a = 64'h21EFFFFFFFFFFFFF; assign b = 64'h1ADFFFFFFFFFFFFF;

    #10 $display("\n2**-480 * 2**-595:");
    #10 assign a = 64'h21F0000000000000; assign b = 64'h1AC0000000000000;
    #10 assign a = 64'h21FFFFFFFFFFFFFF; assign b = 64'h1ACFFFFFFFFFFFFF;

    #10 $display("\n2**-479 * 2**-596:");
    #10 assign a = 64'h2200000000000000; assign b = 64'h1AB0000000000000;
    #10 assign a = 64'h220FFFFFFFFFFFFF; assign b = 64'h1ABFFFFFFFFFFFFF;

    #10 $display("\n2**-478 * 2**-597:");
    #10 assign a = 64'h2210000000000000; assign b = 64'h1AA0000000000000;
    #10 assign a = 64'h221FFFFFFFFFFFFF; assign b = 64'h1AAFFFFFFFFFFFFF;

    #10 $display("\n2**-477 * 2**-598:");
    #10 assign a = 64'h2220000000000000; assign b = 64'h1A90000000000000;
    #10 assign a = 64'h222FFFFFFFFFFFFF; assign b = 64'h1A9FFFFFFFFFFFFF;

    #10 $display("\n2**-476 * 2**-599:");
    #10 assign a = 64'h2230000000000000; assign b = 64'h1A80000000000000;
    #10 assign a = 64'h223FFFFFFFFFFFFF; assign b = 64'h1A8FFFFFFFFFFFFF;

    #10 $display("\n2**-475 * 2**-600:");
    #10 assign a = 64'h2240000000000000; assign b = 64'h1A70000000000000;
    #10 assign a = 64'h224FFFFFFFFFFFFF; assign b = 64'h1A7FFFFFFFFFFFFF;

    #10 $display("\n2**-474 * 2**-601:");
    #10 assign a = 64'h2250000000000000; assign b = 64'h1A60000000000000;
    #10 assign a = 64'h225FFFFFFFFFFFFF; assign b = 64'h1A6FFFFFFFFFFFFF;

    #10 $display("\n2**-473 * 2**-602:");
    #10 assign a = 64'h2260000000000000; assign b = 64'h1A50000000000000;
    #10 assign a = 64'h226FFFFFFFFFFFFF; assign b = 64'h1A5FFFFFFFFFFFFF;

    #10 $display("\n2**-472 * 2**-603:");
    #10 assign a = 64'h2270000000000000; assign b = 64'h1A40000000000000;
    #10 assign a = 64'h227FFFFFFFFFFFFF; assign b = 64'h1A4FFFFFFFFFFFFF;

    #10 $display("\n2**-471 * 2**-604:");
    #10 assign a = 64'h2280000000000000; assign b = 64'h1A30000000000000;
    #10 assign a = 64'h228FFFFFFFFFFFFF; assign b = 64'h1A3FFFFFFFFFFFFF;

    #10 $display("\n2**-470 * 2**-605:");
    #10 assign a = 64'h2290000000000000; assign b = 64'h1A20000000000000;
    #10 assign a = 64'h229FFFFFFFFFFFFF; assign b = 64'h1A2FFFFFFFFFFFFF;

    #10 $display("\n2**-469 * 2**-606:");
    #10 assign a = 64'h22A0000000000000; assign b = 64'h1A10000000000000;
    #10 assign a = 64'h22AFFFFFFFFFFFFF; assign b = 64'h1A1FFFFFFFFFFFFF;

    #10 $display("\n2**-468 * 2**-607:");
    #10 assign a = 64'h22B0000000000000; assign b = 64'h1A00000000000000;
    #10 assign a = 64'h22BFFFFFFFFFFFFF; assign b = 64'h1A0FFFFFFFFFFFFF;

    #10 $display("\n2**-467 * 2**-608:");
    #10 assign a = 64'h22C0000000000000; assign b = 64'h19F0000000000000;
    #10 assign a = 64'h22CFFFFFFFFFFFFF; assign b = 64'h19FFFFFFFFFFFFFF;

    #10 $display("\n2**-466 * 2**-609:");
    #10 assign a = 64'h22D0000000000000; assign b = 64'h19E0000000000000;
    #10 assign a = 64'h22DFFFFFFFFFFFFF; assign b = 64'h19EFFFFFFFFFFFFF;

    #10 $display("\n2**-465 * 2**-610:");
    #10 assign a = 64'h22E0000000000000; assign b = 64'h19D0000000000000;
    #10 assign a = 64'h22EFFFFFFFFFFFFF; assign b = 64'h19DFFFFFFFFFFFFF;

    #10 $display("\n2**-464 * 2**-611:");
    #10 assign a = 64'h22F0000000000000; assign b = 64'h19C0000000000000;
    #10 assign a = 64'h22FFFFFFFFFFFFFF; assign b = 64'h19CFFFFFFFFFFFFF;

    #10 $display("\n2**-463 * 2**-612:");
    #10 assign a = 64'h2300000000000000; assign b = 64'h19B0000000000000;
    #10 assign a = 64'h230FFFFFFFFFFFFF; assign b = 64'h19BFFFFFFFFFFFFF;

    #10 $display("\n2**-462 * 2**-613:");
    #10 assign a = 64'h2310000000000000; assign b = 64'h19A0000000000000;
    #10 assign a = 64'h231FFFFFFFFFFFFF; assign b = 64'h19AFFFFFFFFFFFFF;

    #10 $display("\n2**-461 * 2**-614:");
    #10 assign a = 64'h2320000000000000; assign b = 64'h1990000000000000;
    #10 assign a = 64'h232FFFFFFFFFFFFF; assign b = 64'h199FFFFFFFFFFFFF;

    #10 $display("\n2**-460 * 2**-615:");
    #10 assign a = 64'h2330000000000000; assign b = 64'h1980000000000000;
    #10 assign a = 64'h233FFFFFFFFFFFFF; assign b = 64'h198FFFFFFFFFFFFF;

    #10 $display("\n2**-459 * 2**-616:");
    #10 assign a = 64'h2340000000000000; assign b = 64'h1970000000000000;
    #10 assign a = 64'h234FFFFFFFFFFFFF; assign b = 64'h197FFFFFFFFFFFFF;

    #10 $display("\n2**-458 * 2**-617:");
    #10 assign a = 64'h2350000000000000; assign b = 64'h1960000000000000;
    #10 assign a = 64'h235FFFFFFFFFFFFF; assign b = 64'h196FFFFFFFFFFFFF;

    #10 $display("\n2**-457 * 2**-618:");
    #10 assign a = 64'h2360000000000000; assign b = 64'h1950000000000000;
    #10 assign a = 64'h236FFFFFFFFFFFFF; assign b = 64'h195FFFFFFFFFFFFF;

    #10 $display("\n2**-456 * 2**-619:");
    #10 assign a = 64'h2370000000000000; assign b = 64'h1940000000000000;
    #10 assign a = 64'h237FFFFFFFFFFFFF; assign b = 64'h194FFFFFFFFFFFFF;

    #10 $display("\n2**-455 * 2**-620:");
    #10 assign a = 64'h2380000000000000; assign b = 64'h1930000000000000;
    #10 assign a = 64'h238FFFFFFFFFFFFF; assign b = 64'h193FFFFFFFFFFFFF;

    #10 $display("\n2**-454 * 2**-621:");
    #10 assign a = 64'h2390000000000000; assign b = 64'h1920000000000000;
    #10 assign a = 64'h239FFFFFFFFFFFFF; assign b = 64'h192FFFFFFFFFFFFF;

    #10 $display("\n2**-453 * 2**-622:");
    #10 assign a = 64'h23A0000000000000; assign b = 64'h1910000000000000;
    #10 assign a = 64'h23AFFFFFFFFFFFFF; assign b = 64'h191FFFFFFFFFFFFF;

    #10 $display("\n2**-452 * 2**-623:");
    #10 assign a = 64'h23B0000000000000; assign b = 64'h1900000000000000;
    #10 assign a = 64'h23BFFFFFFFFFFFFF; assign b = 64'h190FFFFFFFFFFFFF;

    #10 $display("\n2**-451 * 2**-624:");
    #10 assign a = 64'h23C0000000000000; assign b = 64'h18F0000000000000;
    #10 assign a = 64'h23CFFFFFFFFFFFFF; assign b = 64'h18FFFFFFFFFFFFFF;

    #10 $display("\n2**-450 * 2**-625:");
    #10 assign a = 64'h23D0000000000000; assign b = 64'h18E0000000000000;
    #10 assign a = 64'h23DFFFFFFFFFFFFF; assign b = 64'h18EFFFFFFFFFFFFF;

    #10 $display("\n2**-449 * 2**-626:");
    #10 assign a = 64'h23E0000000000000; assign b = 64'h18D0000000000000;
    #10 assign a = 64'h23EFFFFFFFFFFFFF; assign b = 64'h18DFFFFFFFFFFFFF;

    #10 $display("\n2**-448 * 2**-627:");
    #10 assign a = 64'h23F0000000000000; assign b = 64'h18C0000000000000;
    #10 assign a = 64'h23FFFFFFFFFFFFFF; assign b = 64'h18CFFFFFFFFFFFFF;

    #10 $display("\n2**-447 * 2**-628:");
    #10 assign a = 64'h2400000000000000; assign b = 64'h18B0000000000000;
    #10 assign a = 64'h240FFFFFFFFFFFFF; assign b = 64'h18BFFFFFFFFFFFFF;

    #10 $display("\n2**-446 * 2**-629:");
    #10 assign a = 64'h2410000000000000; assign b = 64'h18A0000000000000;
    #10 assign a = 64'h241FFFFFFFFFFFFF; assign b = 64'h18AFFFFFFFFFFFFF;

    #10 $display("\n2**-445 * 2**-630:");
    #10 assign a = 64'h2420000000000000; assign b = 64'h1890000000000000;
    #10 assign a = 64'h242FFFFFFFFFFFFF; assign b = 64'h189FFFFFFFFFFFFF;

    #10 $display("\n2**-444 * 2**-631:");
    #10 assign a = 64'h2430000000000000; assign b = 64'h1880000000000000;
    #10 assign a = 64'h243FFFFFFFFFFFFF; assign b = 64'h188FFFFFFFFFFFFF;

    #10 $display("\n2**-443 * 2**-632:");
    #10 assign a = 64'h2440000000000000; assign b = 64'h1870000000000000;
    #10 assign a = 64'h244FFFFFFFFFFFFF; assign b = 64'h187FFFFFFFFFFFFF;

    #10 $display("\n2**-442 * 2**-633:");
    #10 assign a = 64'h2450000000000000; assign b = 64'h1860000000000000;
    #10 assign a = 64'h245FFFFFFFFFFFFF; assign b = 64'h186FFFFFFFFFFFFF;

    #10 $display("\n2**-441 * 2**-634:");
    #10 assign a = 64'h2460000000000000; assign b = 64'h1850000000000000;
    #10 assign a = 64'h246FFFFFFFFFFFFF; assign b = 64'h185FFFFFFFFFFFFF;

    #10 $display("\n2**-440 * 2**-635:");
    #10 assign a = 64'h2470000000000000; assign b = 64'h1840000000000000;
    #10 assign a = 64'h247FFFFFFFFFFFFF; assign b = 64'h184FFFFFFFFFFFFF;

    #10 $display("\n2**-439 * 2**-636:");
    #10 assign a = 64'h2480000000000000; assign b = 64'h1830000000000000;
    #10 assign a = 64'h248FFFFFFFFFFFFF; assign b = 64'h183FFFFFFFFFFFFF;

    #10 $display("\n2**-438 * 2**-637:");
    #10 assign a = 64'h2490000000000000; assign b = 64'h1820000000000000;
    #10 assign a = 64'h249FFFFFFFFFFFFF; assign b = 64'h182FFFFFFFFFFFFF;

    #10 $display("\n2**-437 * 2**-638:");
    #10 assign a = 64'h24A0000000000000; assign b = 64'h1810000000000000;
    #10 assign a = 64'h24AFFFFFFFFFFFFF; assign b = 64'h181FFFFFFFFFFFFF;

    #10 $display("\n2**-436 * 2**-639:");
    #10 assign a = 64'h24B0000000000000; assign b = 64'h1800000000000000;
    #10 assign a = 64'h24BFFFFFFFFFFFFF; assign b = 64'h180FFFFFFFFFFFFF;

    #10 $display("\n2**-435 * 2**-640:");
    #10 assign a = 64'h24C0000000000000; assign b = 64'h17F0000000000000;
    #10 assign a = 64'h24CFFFFFFFFFFFFF; assign b = 64'h17FFFFFFFFFFFFFF;

    #10 $display("\n2**-434 * 2**-641:");
    #10 assign a = 64'h24D0000000000000; assign b = 64'h17E0000000000000;
    #10 assign a = 64'h24DFFFFFFFFFFFFF; assign b = 64'h17EFFFFFFFFFFFFF;

    #10 $display("\n2**-433 * 2**-642:");
    #10 assign a = 64'h24E0000000000000; assign b = 64'h17D0000000000000;
    #10 assign a = 64'h24EFFFFFFFFFFFFF; assign b = 64'h17DFFFFFFFFFFFFF;

    #10 $display("\n2**-432 * 2**-643:");
    #10 assign a = 64'h24F0000000000000; assign b = 64'h17C0000000000000;
    #10 assign a = 64'h24FFFFFFFFFFFFFF; assign b = 64'h17CFFFFFFFFFFFFF;

    #10 $display("\n2**-431 * 2**-644:");
    #10 assign a = 64'h2500000000000000; assign b = 64'h17B0000000000000;
    #10 assign a = 64'h250FFFFFFFFFFFFF; assign b = 64'h17BFFFFFFFFFFFFF;

    #10 $display("\n2**-430 * 2**-645:");
    #10 assign a = 64'h2510000000000000; assign b = 64'h17A0000000000000;
    #10 assign a = 64'h251FFFFFFFFFFFFF; assign b = 64'h17AFFFFFFFFFFFFF;

    #10 $display("\n2**-429 * 2**-646:");
    #10 assign a = 64'h2520000000000000; assign b = 64'h1790000000000000;
    #10 assign a = 64'h252FFFFFFFFFFFFF; assign b = 64'h179FFFFFFFFFFFFF;

    #10 $display("\n2**-428 * 2**-647:");
    #10 assign a = 64'h2530000000000000; assign b = 64'h1780000000000000;
    #10 assign a = 64'h253FFFFFFFFFFFFF; assign b = 64'h178FFFFFFFFFFFFF;

    #10 $display("\n2**-427 * 2**-648:");
    #10 assign a = 64'h2540000000000000; assign b = 64'h1770000000000000;
    #10 assign a = 64'h254FFFFFFFFFFFFF; assign b = 64'h177FFFFFFFFFFFFF;

    #10 $display("\n2**-426 * 2**-649:");
    #10 assign a = 64'h2550000000000000; assign b = 64'h1760000000000000;
    #10 assign a = 64'h255FFFFFFFFFFFFF; assign b = 64'h176FFFFFFFFFFFFF;

    #10 $display("\n2**-425 * 2**-650:");
    #10 assign a = 64'h2560000000000000; assign b = 64'h1750000000000000;
    #10 assign a = 64'h256FFFFFFFFFFFFF; assign b = 64'h175FFFFFFFFFFFFF;

    #10 $display("\n2**-424 * 2**-651:");
    #10 assign a = 64'h2570000000000000; assign b = 64'h1740000000000000;
    #10 assign a = 64'h257FFFFFFFFFFFFF; assign b = 64'h174FFFFFFFFFFFFF;

    #10 $display("\n2**-423 * 2**-652:");
    #10 assign a = 64'h2580000000000000; assign b = 64'h1730000000000000;
    #10 assign a = 64'h258FFFFFFFFFFFFF; assign b = 64'h173FFFFFFFFFFFFF;

    #10 $display("\n2**-422 * 2**-653:");
    #10 assign a = 64'h2590000000000000; assign b = 64'h1720000000000000;
    #10 assign a = 64'h259FFFFFFFFFFFFF; assign b = 64'h172FFFFFFFFFFFFF;

    #10 $display("\n2**-421 * 2**-654:");
    #10 assign a = 64'h25A0000000000000; assign b = 64'h1710000000000000;
    #10 assign a = 64'h25AFFFFFFFFFFFFF; assign b = 64'h171FFFFFFFFFFFFF;

    #10 $display("\n2**-420 * 2**-655:");
    #10 assign a = 64'h25B0000000000000; assign b = 64'h1700000000000000;
    #10 assign a = 64'h25BFFFFFFFFFFFFF; assign b = 64'h170FFFFFFFFFFFFF;

    #10 $display("\n2**-419 * 2**-656:");
    #10 assign a = 64'h25C0000000000000; assign b = 64'h16F0000000000000;
    #10 assign a = 64'h25CFFFFFFFFFFFFF; assign b = 64'h16FFFFFFFFFFFFFF;

    #10 $display("\n2**-418 * 2**-657:");
    #10 assign a = 64'h25D0000000000000; assign b = 64'h16E0000000000000;
    #10 assign a = 64'h25DFFFFFFFFFFFFF; assign b = 64'h16EFFFFFFFFFFFFF;

    #10 $display("\n2**-417 * 2**-658:");
    #10 assign a = 64'h25E0000000000000; assign b = 64'h16D0000000000000;
    #10 assign a = 64'h25EFFFFFFFFFFFFF; assign b = 64'h16DFFFFFFFFFFFFF;

    #10 $display("\n2**-416 * 2**-659:");
    #10 assign a = 64'h25F0000000000000; assign b = 64'h16C0000000000000;
    #10 assign a = 64'h25FFFFFFFFFFFFFF; assign b = 64'h16CFFFFFFFFFFFFF;

    #10 $display("\n2**-415 * 2**-660:");
    #10 assign a = 64'h2600000000000000; assign b = 64'h16B0000000000000;
    #10 assign a = 64'h260FFFFFFFFFFFFF; assign b = 64'h16BFFFFFFFFFFFFF;

    #10 $display("\n2**-414 * 2**-661:");
    #10 assign a = 64'h2610000000000000; assign b = 64'h16A0000000000000;
    #10 assign a = 64'h261FFFFFFFFFFFFF; assign b = 64'h16AFFFFFFFFFFFFF;

    #10 $display("\n2**-413 * 2**-662:");
    #10 assign a = 64'h2620000000000000; assign b = 64'h1690000000000000;
    #10 assign a = 64'h262FFFFFFFFFFFFF; assign b = 64'h169FFFFFFFFFFFFF;

    #10 $display("\n2**-412 * 2**-663:");
    #10 assign a = 64'h2630000000000000; assign b = 64'h1680000000000000;
    #10 assign a = 64'h263FFFFFFFFFFFFF; assign b = 64'h168FFFFFFFFFFFFF;

    #10 $display("\n2**-411 * 2**-664:");
    #10 assign a = 64'h2640000000000000; assign b = 64'h1670000000000000;
    #10 assign a = 64'h264FFFFFFFFFFFFF; assign b = 64'h167FFFFFFFFFFFFF;

    #10 $display("\n2**-410 * 2**-665:");
    #10 assign a = 64'h2650000000000000; assign b = 64'h1660000000000000;
    #10 assign a = 64'h265FFFFFFFFFFFFF; assign b = 64'h166FFFFFFFFFFFFF;

    #10 $display("\n2**-409 * 2**-666:");
    #10 assign a = 64'h2660000000000000; assign b = 64'h1650000000000000;
    #10 assign a = 64'h266FFFFFFFFFFFFF; assign b = 64'h165FFFFFFFFFFFFF;

    #10 $display("\n2**-408 * 2**-667:");
    #10 assign a = 64'h2670000000000000; assign b = 64'h1640000000000000;
    #10 assign a = 64'h267FFFFFFFFFFFFF; assign b = 64'h164FFFFFFFFFFFFF;

    #10 $display("\n2**-407 * 2**-668:");
    #10 assign a = 64'h2680000000000000; assign b = 64'h1630000000000000;
    #10 assign a = 64'h268FFFFFFFFFFFFF; assign b = 64'h163FFFFFFFFFFFFF;

    #10 $display("\n2**-406 * 2**-669:");
    #10 assign a = 64'h2690000000000000; assign b = 64'h1620000000000000;
    #10 assign a = 64'h269FFFFFFFFFFFFF; assign b = 64'h162FFFFFFFFFFFFF;

    #10 $display("\n2**-405 * 2**-670:");
    #10 assign a = 64'h26A0000000000000; assign b = 64'h1610000000000000;
    #10 assign a = 64'h26AFFFFFFFFFFFFF; assign b = 64'h161FFFFFFFFFFFFF;

    #10 $display("\n2**-404 * 2**-671:");
    #10 assign a = 64'h26B0000000000000; assign b = 64'h1600000000000000;
    #10 assign a = 64'h26BFFFFFFFFFFFFF; assign b = 64'h160FFFFFFFFFFFFF;

    #10 $display("\n2**-403 * 2**-672:");
    #10 assign a = 64'h26C0000000000000; assign b = 64'h15F0000000000000;
    #10 assign a = 64'h26CFFFFFFFFFFFFF; assign b = 64'h15FFFFFFFFFFFFFF;

    #10 $display("\n2**-402 * 2**-673:");
    #10 assign a = 64'h26D0000000000000; assign b = 64'h15E0000000000000;
    #10 assign a = 64'h26DFFFFFFFFFFFFF; assign b = 64'h15EFFFFFFFFFFFFF;

    #10 $display("\n2**-401 * 2**-674:");
    #10 assign a = 64'h26E0000000000000; assign b = 64'h15D0000000000000;
    #10 assign a = 64'h26EFFFFFFFFFFFFF; assign b = 64'h15DFFFFFFFFFFFFF;

    #10 $display("\n2**-400 * 2**-675:");
    #10 assign a = 64'h26F0000000000000; assign b = 64'h15C0000000000000;
    #10 assign a = 64'h26FFFFFFFFFFFFFF; assign b = 64'h15CFFFFFFFFFFFFF;

    #10 $display("\n2**-399 * 2**-676:");
    #10 assign a = 64'h2700000000000000; assign b = 64'h15B0000000000000;
    #10 assign a = 64'h270FFFFFFFFFFFFF; assign b = 64'h15BFFFFFFFFFFFFF;

    #10 $display("\n2**-398 * 2**-677:");
    #10 assign a = 64'h2710000000000000; assign b = 64'h15A0000000000000;
    #10 assign a = 64'h271FFFFFFFFFFFFF; assign b = 64'h15AFFFFFFFFFFFFF;

    #10 $display("\n2**-397 * 2**-678:");
    #10 assign a = 64'h2720000000000000; assign b = 64'h1590000000000000;
    #10 assign a = 64'h272FFFFFFFFFFFFF; assign b = 64'h159FFFFFFFFFFFFF;

    #10 $display("\n2**-396 * 2**-679:");
    #10 assign a = 64'h2730000000000000; assign b = 64'h1580000000000000;
    #10 assign a = 64'h273FFFFFFFFFFFFF; assign b = 64'h158FFFFFFFFFFFFF;

    #10 $display("\n2**-395 * 2**-680:");
    #10 assign a = 64'h2740000000000000; assign b = 64'h1570000000000000;
    #10 assign a = 64'h274FFFFFFFFFFFFF; assign b = 64'h157FFFFFFFFFFFFF;

    #10 $display("\n2**-394 * 2**-681:");
    #10 assign a = 64'h2750000000000000; assign b = 64'h1560000000000000;
    #10 assign a = 64'h275FFFFFFFFFFFFF; assign b = 64'h156FFFFFFFFFFFFF;

    #10 $display("\n2**-393 * 2**-682:");
    #10 assign a = 64'h2760000000000000; assign b = 64'h1550000000000000;
    #10 assign a = 64'h276FFFFFFFFFFFFF; assign b = 64'h155FFFFFFFFFFFFF;

    #10 $display("\n2**-392 * 2**-683:");
    #10 assign a = 64'h2770000000000000; assign b = 64'h1540000000000000;
    #10 assign a = 64'h277FFFFFFFFFFFFF; assign b = 64'h154FFFFFFFFFFFFF;

    #10 $display("\n2**-391 * 2**-684:");
    #10 assign a = 64'h2780000000000000; assign b = 64'h1530000000000000;
    #10 assign a = 64'h278FFFFFFFFFFFFF; assign b = 64'h153FFFFFFFFFFFFF;

    #10 $display("\n2**-390 * 2**-685:");
    #10 assign a = 64'h2790000000000000; assign b = 64'h1520000000000000;
    #10 assign a = 64'h279FFFFFFFFFFFFF; assign b = 64'h152FFFFFFFFFFFFF;

    #10 $display("\n2**-389 * 2**-686:");
    #10 assign a = 64'h27A0000000000000; assign b = 64'h1510000000000000;
    #10 assign a = 64'h27AFFFFFFFFFFFFF; assign b = 64'h151FFFFFFFFFFFFF;

    #10 $display("\n2**-388 * 2**-687:");
    #10 assign a = 64'h27B0000000000000; assign b = 64'h1500000000000000;
    #10 assign a = 64'h27BFFFFFFFFFFFFF; assign b = 64'h150FFFFFFFFFFFFF;

    #10 $display("\n2**-387 * 2**-688:");
    #10 assign a = 64'h27C0000000000000; assign b = 64'h14F0000000000000;
    #10 assign a = 64'h27CFFFFFFFFFFFFF; assign b = 64'h14FFFFFFFFFFFFFF;

    #10 $display("\n2**-386 * 2**-689:");
    #10 assign a = 64'h27D0000000000000; assign b = 64'h14E0000000000000;
    #10 assign a = 64'h27DFFFFFFFFFFFFF; assign b = 64'h14EFFFFFFFFFFFFF;

    #10 $display("\n2**-385 * 2**-690:");
    #10 assign a = 64'h27E0000000000000; assign b = 64'h14D0000000000000;
    #10 assign a = 64'h27EFFFFFFFFFFFFF; assign b = 64'h14DFFFFFFFFFFFFF;

    #10 $display("\n2**-384 * 2**-691:");
    #10 assign a = 64'h27F0000000000000; assign b = 64'h14C0000000000000;
    #10 assign a = 64'h27FFFFFFFFFFFFFF; assign b = 64'h14CFFFFFFFFFFFFF;

    #10 $display("\n2**-383 * 2**-692:");
    #10 assign a = 64'h2800000000000000; assign b = 64'h14B0000000000000;
    #10 assign a = 64'h280FFFFFFFFFFFFF; assign b = 64'h14BFFFFFFFFFFFFF;

    #10 $display("\n2**-382 * 2**-693:");
    #10 assign a = 64'h2810000000000000; assign b = 64'h14A0000000000000;
    #10 assign a = 64'h281FFFFFFFFFFFFF; assign b = 64'h14AFFFFFFFFFFFFF;

    #10 $display("\n2**-381 * 2**-694:");
    #10 assign a = 64'h2820000000000000; assign b = 64'h1490000000000000;
    #10 assign a = 64'h282FFFFFFFFFFFFF; assign b = 64'h149FFFFFFFFFFFFF;

    #10 $display("\n2**-380 * 2**-695:");
    #10 assign a = 64'h2830000000000000; assign b = 64'h1480000000000000;
    #10 assign a = 64'h283FFFFFFFFFFFFF; assign b = 64'h148FFFFFFFFFFFFF;

    #10 $display("\n2**-379 * 2**-696:");
    #10 assign a = 64'h2840000000000000; assign b = 64'h1470000000000000;
    #10 assign a = 64'h284FFFFFFFFFFFFF; assign b = 64'h147FFFFFFFFFFFFF;

    #10 $display("\n2**-378 * 2**-697:");
    #10 assign a = 64'h2850000000000000; assign b = 64'h1460000000000000;
    #10 assign a = 64'h285FFFFFFFFFFFFF; assign b = 64'h146FFFFFFFFFFFFF;

    #10 $display("\n2**-377 * 2**-698:");
    #10 assign a = 64'h2860000000000000; assign b = 64'h1450000000000000;
    #10 assign a = 64'h286FFFFFFFFFFFFF; assign b = 64'h145FFFFFFFFFFFFF;

    #10 $display("\n2**-376 * 2**-699:");
    #10 assign a = 64'h2870000000000000; assign b = 64'h1440000000000000;
    #10 assign a = 64'h287FFFFFFFFFFFFF; assign b = 64'h144FFFFFFFFFFFFF;

    #10 $display("\n2**-375 * 2**-700:");
    #10 assign a = 64'h2880000000000000; assign b = 64'h1430000000000000;
    #10 assign a = 64'h288FFFFFFFFFFFFF; assign b = 64'h143FFFFFFFFFFFFF;

    #10 $display("\n2**-374 * 2**-701:");
    #10 assign a = 64'h2890000000000000; assign b = 64'h1420000000000000;
    #10 assign a = 64'h289FFFFFFFFFFFFF; assign b = 64'h142FFFFFFFFFFFFF;

    #10 $display("\n2**-373 * 2**-702:");
    #10 assign a = 64'h28A0000000000000; assign b = 64'h1410000000000000;
    #10 assign a = 64'h28AFFFFFFFFFFFFF; assign b = 64'h141FFFFFFFFFFFFF;

    #10 $display("\n2**-372 * 2**-703:");
    #10 assign a = 64'h28B0000000000000; assign b = 64'h1400000000000000;
    #10 assign a = 64'h28BFFFFFFFFFFFFF; assign b = 64'h140FFFFFFFFFFFFF;

    #10 $display("\n2**-371 * 2**-704:");
    #10 assign a = 64'h28C0000000000000; assign b = 64'h13F0000000000000;
    #10 assign a = 64'h28CFFFFFFFFFFFFF; assign b = 64'h13FFFFFFFFFFFFFF;

    #10 $display("\n2**-370 * 2**-705:");
    #10 assign a = 64'h28D0000000000000; assign b = 64'h13E0000000000000;
    #10 assign a = 64'h28DFFFFFFFFFFFFF; assign b = 64'h13EFFFFFFFFFFFFF;

    #10 $display("\n2**-369 * 2**-706:");
    #10 assign a = 64'h28E0000000000000; assign b = 64'h13D0000000000000;
    #10 assign a = 64'h28EFFFFFFFFFFFFF; assign b = 64'h13DFFFFFFFFFFFFF;

    #10 $display("\n2**-368 * 2**-707:");
    #10 assign a = 64'h28F0000000000000; assign b = 64'h13C0000000000000;
    #10 assign a = 64'h28FFFFFFFFFFFFFF; assign b = 64'h13CFFFFFFFFFFFFF;

    #10 $display("\n2**-367 * 2**-708:");
    #10 assign a = 64'h2900000000000000; assign b = 64'h13B0000000000000;
    #10 assign a = 64'h290FFFFFFFFFFFFF; assign b = 64'h13BFFFFFFFFFFFFF;

    #10 $display("\n2**-366 * 2**-709:");
    #10 assign a = 64'h2910000000000000; assign b = 64'h13A0000000000000;
    #10 assign a = 64'h291FFFFFFFFFFFFF; assign b = 64'h13AFFFFFFFFFFFFF;

    #10 $display("\n2**-365 * 2**-710:");
    #10 assign a = 64'h2920000000000000; assign b = 64'h1390000000000000;
    #10 assign a = 64'h292FFFFFFFFFFFFF; assign b = 64'h139FFFFFFFFFFFFF;

    #10 $display("\n2**-364 * 2**-711:");
    #10 assign a = 64'h2930000000000000; assign b = 64'h1380000000000000;
    #10 assign a = 64'h293FFFFFFFFFFFFF; assign b = 64'h138FFFFFFFFFFFFF;

    #10 $display("\n2**-363 * 2**-712:");
    #10 assign a = 64'h2940000000000000; assign b = 64'h1370000000000000;
    #10 assign a = 64'h294FFFFFFFFFFFFF; assign b = 64'h137FFFFFFFFFFFFF;

    #10 $display("\n2**-362 * 2**-713:");
    #10 assign a = 64'h2950000000000000; assign b = 64'h1360000000000000;
    #10 assign a = 64'h295FFFFFFFFFFFFF; assign b = 64'h136FFFFFFFFFFFFF;

    #10 $display("\n2**-361 * 2**-714:");
    #10 assign a = 64'h2960000000000000; assign b = 64'h1350000000000000;
    #10 assign a = 64'h296FFFFFFFFFFFFF; assign b = 64'h135FFFFFFFFFFFFF;

    #10 $display("\n2**-360 * 2**-715:");
    #10 assign a = 64'h2970000000000000; assign b = 64'h1340000000000000;
    #10 assign a = 64'h297FFFFFFFFFFFFF; assign b = 64'h134FFFFFFFFFFFFF;

    #10 $display("\n2**-359 * 2**-716:");
    #10 assign a = 64'h2980000000000000; assign b = 64'h1330000000000000;
    #10 assign a = 64'h298FFFFFFFFFFFFF; assign b = 64'h133FFFFFFFFFFFFF;

    #10 $display("\n2**-358 * 2**-717:");
    #10 assign a = 64'h2990000000000000; assign b = 64'h1320000000000000;
    #10 assign a = 64'h299FFFFFFFFFFFFF; assign b = 64'h132FFFFFFFFFFFFF;

    #10 $display("\n2**-357 * 2**-718:");
    #10 assign a = 64'h29A0000000000000; assign b = 64'h1310000000000000;
    #10 assign a = 64'h29AFFFFFFFFFFFFF; assign b = 64'h131FFFFFFFFFFFFF;

    #10 $display("\n2**-356 * 2**-719:");
    #10 assign a = 64'h29B0000000000000; assign b = 64'h1300000000000000;
    #10 assign a = 64'h29BFFFFFFFFFFFFF; assign b = 64'h130FFFFFFFFFFFFF;

    #10 $display("\n2**-355 * 2**-720:");
    #10 assign a = 64'h29C0000000000000; assign b = 64'h12F0000000000000;
    #10 assign a = 64'h29CFFFFFFFFFFFFF; assign b = 64'h12FFFFFFFFFFFFFF;

    #10 $display("\n2**-354 * 2**-721:");
    #10 assign a = 64'h29D0000000000000; assign b = 64'h12E0000000000000;
    #10 assign a = 64'h29DFFFFFFFFFFFFF; assign b = 64'h12EFFFFFFFFFFFFF;

    #10 $display("\n2**-353 * 2**-722:");
    #10 assign a = 64'h29E0000000000000; assign b = 64'h12D0000000000000;
    #10 assign a = 64'h29EFFFFFFFFFFFFF; assign b = 64'h12DFFFFFFFFFFFFF;

    #10 $display("\n2**-352 * 2**-723:");
    #10 assign a = 64'h29F0000000000000; assign b = 64'h12C0000000000000;
    #10 assign a = 64'h29FFFFFFFFFFFFFF; assign b = 64'h12CFFFFFFFFFFFFF;

    #10 $display("\n2**-351 * 2**-724:");
    #10 assign a = 64'h2A00000000000000; assign b = 64'h12B0000000000000;
    #10 assign a = 64'h2A0FFFFFFFFFFFFF; assign b = 64'h12BFFFFFFFFFFFFF;

    #10 $display("\n2**-350 * 2**-725:");
    #10 assign a = 64'h2A10000000000000; assign b = 64'h12A0000000000000;
    #10 assign a = 64'h2A1FFFFFFFFFFFFF; assign b = 64'h12AFFFFFFFFFFFFF;

    #10 $display("\n2**-349 * 2**-726:");
    #10 assign a = 64'h2A20000000000000; assign b = 64'h1290000000000000;
    #10 assign a = 64'h2A2FFFFFFFFFFFFF; assign b = 64'h129FFFFFFFFFFFFF;

    #10 $display("\n2**-348 * 2**-727:");
    #10 assign a = 64'h2A30000000000000; assign b = 64'h1280000000000000;
    #10 assign a = 64'h2A3FFFFFFFFFFFFF; assign b = 64'h128FFFFFFFFFFFFF;

    #10 $display("\n2**-347 * 2**-728:");
    #10 assign a = 64'h2A40000000000000; assign b = 64'h1270000000000000;
    #10 assign a = 64'h2A4FFFFFFFFFFFFF; assign b = 64'h127FFFFFFFFFFFFF;

    #10 $display("\n2**-346 * 2**-729:");
    #10 assign a = 64'h2A50000000000000; assign b = 64'h1260000000000000;
    #10 assign a = 64'h2A5FFFFFFFFFFFFF; assign b = 64'h126FFFFFFFFFFFFF;

    #10 $display("\n2**-345 * 2**-730:");
    #10 assign a = 64'h2A60000000000000; assign b = 64'h1250000000000000;
    #10 assign a = 64'h2A6FFFFFFFFFFFFF; assign b = 64'h125FFFFFFFFFFFFF;

    #10 $display("\n2**-344 * 2**-731:");
    #10 assign a = 64'h2A70000000000000; assign b = 64'h1240000000000000;
    #10 assign a = 64'h2A7FFFFFFFFFFFFF; assign b = 64'h124FFFFFFFFFFFFF;

    #10 $display("\n2**-343 * 2**-732:");
    #10 assign a = 64'h2A80000000000000; assign b = 64'h1230000000000000;
    #10 assign a = 64'h2A8FFFFFFFFFFFFF; assign b = 64'h123FFFFFFFFFFFFF;

    #10 $display("\n2**-342 * 2**-733:");
    #10 assign a = 64'h2A90000000000000; assign b = 64'h1220000000000000;
    #10 assign a = 64'h2A9FFFFFFFFFFFFF; assign b = 64'h122FFFFFFFFFFFFF;

    #10 $display("\n2**-341 * 2**-734:");
    #10 assign a = 64'h2AA0000000000000; assign b = 64'h1210000000000000;
    #10 assign a = 64'h2AAFFFFFFFFFFFFF; assign b = 64'h121FFFFFFFFFFFFF;

    #10 $display("\n2**-340 * 2**-735:");
    #10 assign a = 64'h2AB0000000000000; assign b = 64'h1200000000000000;
    #10 assign a = 64'h2ABFFFFFFFFFFFFF; assign b = 64'h120FFFFFFFFFFFFF;

    #10 $display("\n2**-339 * 2**-736:");
    #10 assign a = 64'h2AC0000000000000; assign b = 64'h11F0000000000000;
    #10 assign a = 64'h2ACFFFFFFFFFFFFF; assign b = 64'h11FFFFFFFFFFFFFF;

    #10 $display("\n2**-338 * 2**-737:");
    #10 assign a = 64'h2AD0000000000000; assign b = 64'h11E0000000000000;
    #10 assign a = 64'h2ADFFFFFFFFFFFFF; assign b = 64'h11EFFFFFFFFFFFFF;

    #10 $display("\n2**-337 * 2**-738:");
    #10 assign a = 64'h2AE0000000000000; assign b = 64'h11D0000000000000;
    #10 assign a = 64'h2AEFFFFFFFFFFFFF; assign b = 64'h11DFFFFFFFFFFFFF;

    #10 $display("\n2**-336 * 2**-739:");
    #10 assign a = 64'h2AF0000000000000; assign b = 64'h11C0000000000000;
    #10 assign a = 64'h2AFFFFFFFFFFFFFF; assign b = 64'h11CFFFFFFFFFFFFF;

    #10 $display("\n2**-335 * 2**-740:");
    #10 assign a = 64'h2B00000000000000; assign b = 64'h11B0000000000000;
    #10 assign a = 64'h2B0FFFFFFFFFFFFF; assign b = 64'h11BFFFFFFFFFFFFF;

    #10 $display("\n2**-334 * 2**-741:");
    #10 assign a = 64'h2B10000000000000; assign b = 64'h11A0000000000000;
    #10 assign a = 64'h2B1FFFFFFFFFFFFF; assign b = 64'h11AFFFFFFFFFFFFF;

    #10 $display("\n2**-333 * 2**-742:");
    #10 assign a = 64'h2B20000000000000; assign b = 64'h1190000000000000;
    #10 assign a = 64'h2B2FFFFFFFFFFFFF; assign b = 64'h119FFFFFFFFFFFFF;

    #10 $display("\n2**-332 * 2**-743:");
    #10 assign a = 64'h2B30000000000000; assign b = 64'h1180000000000000;
    #10 assign a = 64'h2B3FFFFFFFFFFFFF; assign b = 64'h118FFFFFFFFFFFFF;

    #10 $display("\n2**-331 * 2**-744:");
    #10 assign a = 64'h2B40000000000000; assign b = 64'h1170000000000000;
    #10 assign a = 64'h2B4FFFFFFFFFFFFF; assign b = 64'h117FFFFFFFFFFFFF;

    #10 $display("\n2**-330 * 2**-745:");
    #10 assign a = 64'h2B50000000000000; assign b = 64'h1160000000000000;
    #10 assign a = 64'h2B5FFFFFFFFFFFFF; assign b = 64'h116FFFFFFFFFFFFF;

    #10 $display("\n2**-329 * 2**-746:");
    #10 assign a = 64'h2B60000000000000; assign b = 64'h1150000000000000;
    #10 assign a = 64'h2B6FFFFFFFFFFFFF; assign b = 64'h115FFFFFFFFFFFFF;

    #10 $display("\n2**-328 * 2**-747:");
    #10 assign a = 64'h2B70000000000000; assign b = 64'h1140000000000000;
    #10 assign a = 64'h2B7FFFFFFFFFFFFF; assign b = 64'h114FFFFFFFFFFFFF;

    #10 $display("\n2**-327 * 2**-748:");
    #10 assign a = 64'h2B80000000000000; assign b = 64'h1130000000000000;
    #10 assign a = 64'h2B8FFFFFFFFFFFFF; assign b = 64'h113FFFFFFFFFFFFF;

    #10 $display("\n2**-326 * 2**-749:");
    #10 assign a = 64'h2B90000000000000; assign b = 64'h1120000000000000;
    #10 assign a = 64'h2B9FFFFFFFFFFFFF; assign b = 64'h112FFFFFFFFFFFFF;

    #10 $display("\n2**-325 * 2**-750:");
    #10 assign a = 64'h2BA0000000000000; assign b = 64'h1110000000000000;
    #10 assign a = 64'h2BAFFFFFFFFFFFFF; assign b = 64'h111FFFFFFFFFFFFF;

    #10 $display("\n2**-324 * 2**-751:");
    #10 assign a = 64'h2BB0000000000000; assign b = 64'h1100000000000000;
    #10 assign a = 64'h2BBFFFFFFFFFFFFF; assign b = 64'h110FFFFFFFFFFFFF;

    #10 $display("\n2**-323 * 2**-752:");
    #10 assign a = 64'h2BC0000000000000; assign b = 64'h10F0000000000000;
    #10 assign a = 64'h2BCFFFFFFFFFFFFF; assign b = 64'h10FFFFFFFFFFFFFF;

    #10 $display("\n2**-322 * 2**-753:");
    #10 assign a = 64'h2BD0000000000000; assign b = 64'h10E0000000000000;
    #10 assign a = 64'h2BDFFFFFFFFFFFFF; assign b = 64'h10EFFFFFFFFFFFFF;

    #10 $display("\n2**-321 * 2**-754:");
    #10 assign a = 64'h2BE0000000000000; assign b = 64'h10D0000000000000;
    #10 assign a = 64'h2BEFFFFFFFFFFFFF; assign b = 64'h10DFFFFFFFFFFFFF;

    #10 $display("\n2**-320 * 2**-755:");
    #10 assign a = 64'h2BF0000000000000; assign b = 64'h10C0000000000000;
    #10 assign a = 64'h2BFFFFFFFFFFFFFF; assign b = 64'h10CFFFFFFFFFFFFF;

    #10 $display("\n2**-319 * 2**-756:");
    #10 assign a = 64'h2C00000000000000; assign b = 64'h10B0000000000000;
    #10 assign a = 64'h2C0FFFFFFFFFFFFF; assign b = 64'h10BFFFFFFFFFFFFF;

    #10 $display("\n2**-318 * 2**-757:");
    #10 assign a = 64'h2C10000000000000; assign b = 64'h10A0000000000000;
    #10 assign a = 64'h2C1FFFFFFFFFFFFF; assign b = 64'h10AFFFFFFFFFFFFF;

    #10 $display("\n2**-317 * 2**-758:");
    #10 assign a = 64'h2C20000000000000; assign b = 64'h1090000000000000;
    #10 assign a = 64'h2C2FFFFFFFFFFFFF; assign b = 64'h109FFFFFFFFFFFFF;

    #10 $display("\n2**-316 * 2**-759:");
    #10 assign a = 64'h2C30000000000000; assign b = 64'h1080000000000000;
    #10 assign a = 64'h2C3FFFFFFFFFFFFF; assign b = 64'h108FFFFFFFFFFFFF;

    #10 $display("\n2**-315 * 2**-760:");
    #10 assign a = 64'h2C40000000000000; assign b = 64'h1070000000000000;
    #10 assign a = 64'h2C4FFFFFFFFFFFFF; assign b = 64'h107FFFFFFFFFFFFF;

    #10 $display("\n2**-314 * 2**-761:");
    #10 assign a = 64'h2C50000000000000; assign b = 64'h1060000000000000;
    #10 assign a = 64'h2C5FFFFFFFFFFFFF; assign b = 64'h106FFFFFFFFFFFFF;

    #10 $display("\n2**-313 * 2**-762:");
    #10 assign a = 64'h2C60000000000000; assign b = 64'h1050000000000000;
    #10 assign a = 64'h2C6FFFFFFFFFFFFF; assign b = 64'h105FFFFFFFFFFFFF;

    #10 $display("\n2**-312 * 2**-763:");
    #10 assign a = 64'h2C70000000000000; assign b = 64'h1040000000000000;
    #10 assign a = 64'h2C7FFFFFFFFFFFFF; assign b = 64'h104FFFFFFFFFFFFF;

    #10 $display("\n2**-311 * 2**-764:");
    #10 assign a = 64'h2C80000000000000; assign b = 64'h1030000000000000;
    #10 assign a = 64'h2C8FFFFFFFFFFFFF; assign b = 64'h103FFFFFFFFFFFFF;

    #10 $display("\n2**-310 * 2**-765:");
    #10 assign a = 64'h2C90000000000000; assign b = 64'h1020000000000000;
    #10 assign a = 64'h2C9FFFFFFFFFFFFF; assign b = 64'h102FFFFFFFFFFFFF;

    #10 $display("\n2**-309 * 2**-766:");
    #10 assign a = 64'h2CA0000000000000; assign b = 64'h1010000000000000;
    #10 assign a = 64'h2CAFFFFFFFFFFFFF; assign b = 64'h101FFFFFFFFFFFFF;

    #10 $display("\n2**-308 * 2**-767:");
    #10 assign a = 64'h2CB0000000000000; assign b = 64'h1000000000000000;
    #10 assign a = 64'h2CBFFFFFFFFFFFFF; assign b = 64'h100FFFFFFFFFFFFF;

    #10 $display("\n2**-307 * 2**-768:");
    #10 assign a = 64'h2CC0000000000000; assign b = 64'h0FF0000000000000;
    #10 assign a = 64'h2CCFFFFFFFFFFFFF; assign b = 64'h0FFFFFFFFFFFFFFF;

    #10 $display("\n2**-306 * 2**-769:");
    #10 assign a = 64'h2CD0000000000000; assign b = 64'h0FE0000000000000;
    #10 assign a = 64'h2CDFFFFFFFFFFFFF; assign b = 64'h0FEFFFFFFFFFFFFF;

    #10 $display("\n2**-305 * 2**-770:");
    #10 assign a = 64'h2CE0000000000000; assign b = 64'h0FD0000000000000;
    #10 assign a = 64'h2CEFFFFFFFFFFFFF; assign b = 64'h0FDFFFFFFFFFFFFF;

    #10 $display("\n2**-304 * 2**-771:");
    #10 assign a = 64'h2CF0000000000000; assign b = 64'h0FC0000000000000;
    #10 assign a = 64'h2CFFFFFFFFFFFFFF; assign b = 64'h0FCFFFFFFFFFFFFF;

    #10 $display("\n2**-303 * 2**-772:");
    #10 assign a = 64'h2D00000000000000; assign b = 64'h0FB0000000000000;
    #10 assign a = 64'h2D0FFFFFFFFFFFFF; assign b = 64'h0FBFFFFFFFFFFFFF;

    #10 $display("\n2**-302 * 2**-773:");
    #10 assign a = 64'h2D10000000000000; assign b = 64'h0FA0000000000000;
    #10 assign a = 64'h2D1FFFFFFFFFFFFF; assign b = 64'h0FAFFFFFFFFFFFFF;

    #10 $display("\n2**-301 * 2**-774:");
    #10 assign a = 64'h2D20000000000000; assign b = 64'h0F90000000000000;
    #10 assign a = 64'h2D2FFFFFFFFFFFFF; assign b = 64'h0F9FFFFFFFFFFFFF;

    #10 $display("\n2**-300 * 2**-775:");
    #10 assign a = 64'h2D30000000000000; assign b = 64'h0F80000000000000;
    #10 assign a = 64'h2D3FFFFFFFFFFFFF; assign b = 64'h0F8FFFFFFFFFFFFF;

    #10 $display("\n2**-299 * 2**-776:");
    #10 assign a = 64'h2D40000000000000; assign b = 64'h0F70000000000000;
    #10 assign a = 64'h2D4FFFFFFFFFFFFF; assign b = 64'h0F7FFFFFFFFFFFFF;

    #10 $display("\n2**-298 * 2**-777:");
    #10 assign a = 64'h2D50000000000000; assign b = 64'h0F60000000000000;
    #10 assign a = 64'h2D5FFFFFFFFFFFFF; assign b = 64'h0F6FFFFFFFFFFFFF;

    #10 $display("\n2**-297 * 2**-778:");
    #10 assign a = 64'h2D60000000000000; assign b = 64'h0F50000000000000;
    #10 assign a = 64'h2D6FFFFFFFFFFFFF; assign b = 64'h0F5FFFFFFFFFFFFF;

    #10 $display("\n2**-296 * 2**-779:");
    #10 assign a = 64'h2D70000000000000; assign b = 64'h0F40000000000000;
    #10 assign a = 64'h2D7FFFFFFFFFFFFF; assign b = 64'h0F4FFFFFFFFFFFFF;

    #10 $display("\n2**-295 * 2**-780:");
    #10 assign a = 64'h2D80000000000000; assign b = 64'h0F30000000000000;
    #10 assign a = 64'h2D8FFFFFFFFFFFFF; assign b = 64'h0F3FFFFFFFFFFFFF;

    #10 $display("\n2**-294 * 2**-781:");
    #10 assign a = 64'h2D90000000000000; assign b = 64'h0F20000000000000;
    #10 assign a = 64'h2D9FFFFFFFFFFFFF; assign b = 64'h0F2FFFFFFFFFFFFF;

    #10 $display("\n2**-293 * 2**-782:");
    #10 assign a = 64'h2DA0000000000000; assign b = 64'h0F10000000000000;
    #10 assign a = 64'h2DAFFFFFFFFFFFFF; assign b = 64'h0F1FFFFFFFFFFFFF;

    #10 $display("\n2**-292 * 2**-783:");
    #10 assign a = 64'h2DB0000000000000; assign b = 64'h0F00000000000000;
    #10 assign a = 64'h2DBFFFFFFFFFFFFF; assign b = 64'h0F0FFFFFFFFFFFFF;

    #10 $display("\n2**-291 * 2**-784:");
    #10 assign a = 64'h2DC0000000000000; assign b = 64'h0EF0000000000000;
    #10 assign a = 64'h2DCFFFFFFFFFFFFF; assign b = 64'h0EFFFFFFFFFFFFFF;

    #10 $display("\n2**-290 * 2**-785:");
    #10 assign a = 64'h2DD0000000000000; assign b = 64'h0EE0000000000000;
    #10 assign a = 64'h2DDFFFFFFFFFFFFF; assign b = 64'h0EEFFFFFFFFFFFFF;

    #10 $display("\n2**-289 * 2**-786:");
    #10 assign a = 64'h2DE0000000000000; assign b = 64'h0ED0000000000000;
    #10 assign a = 64'h2DEFFFFFFFFFFFFF; assign b = 64'h0EDFFFFFFFFFFFFF;

    #10 $display("\n2**-288 * 2**-787:");
    #10 assign a = 64'h2DF0000000000000; assign b = 64'h0EC0000000000000;
    #10 assign a = 64'h2DFFFFFFFFFFFFFF; assign b = 64'h0ECFFFFFFFFFFFFF;

    #10 $display("\n2**-287 * 2**-788:");
    #10 assign a = 64'h2E00000000000000; assign b = 64'h0EB0000000000000;
    #10 assign a = 64'h2E0FFFFFFFFFFFFF; assign b = 64'h0EBFFFFFFFFFFFFF;

    #10 $display("\n2**-286 * 2**-789:");
    #10 assign a = 64'h2E10000000000000; assign b = 64'h0EA0000000000000;
    #10 assign a = 64'h2E1FFFFFFFFFFFFF; assign b = 64'h0EAFFFFFFFFFFFFF;

    #10 $display("\n2**-285 * 2**-790:");
    #10 assign a = 64'h2E20000000000000; assign b = 64'h0E90000000000000;
    #10 assign a = 64'h2E2FFFFFFFFFFFFF; assign b = 64'h0E9FFFFFFFFFFFFF;

    #10 $display("\n2**-284 * 2**-791:");
    #10 assign a = 64'h2E30000000000000; assign b = 64'h0E80000000000000;
    #10 assign a = 64'h2E3FFFFFFFFFFFFF; assign b = 64'h0E8FFFFFFFFFFFFF;

    #10 $display("\n2**-283 * 2**-792:");
    #10 assign a = 64'h2E40000000000000; assign b = 64'h0E70000000000000;
    #10 assign a = 64'h2E4FFFFFFFFFFFFF; assign b = 64'h0E7FFFFFFFFFFFFF;

    #10 $display("\n2**-282 * 2**-793:");
    #10 assign a = 64'h2E50000000000000; assign b = 64'h0E60000000000000;
    #10 assign a = 64'h2E5FFFFFFFFFFFFF; assign b = 64'h0E6FFFFFFFFFFFFF;

    #10 $display("\n2**-281 * 2**-794:");
    #10 assign a = 64'h2E60000000000000; assign b = 64'h0E50000000000000;
    #10 assign a = 64'h2E6FFFFFFFFFFFFF; assign b = 64'h0E5FFFFFFFFFFFFF;

    #10 $display("\n2**-280 * 2**-795:");
    #10 assign a = 64'h2E70000000000000; assign b = 64'h0E40000000000000;
    #10 assign a = 64'h2E7FFFFFFFFFFFFF; assign b = 64'h0E4FFFFFFFFFFFFF;

    #10 $display("\n2**-279 * 2**-796:");
    #10 assign a = 64'h2E80000000000000; assign b = 64'h0E30000000000000;
    #10 assign a = 64'h2E8FFFFFFFFFFFFF; assign b = 64'h0E3FFFFFFFFFFFFF;

    #10 $display("\n2**-278 * 2**-797:");
    #10 assign a = 64'h2E90000000000000; assign b = 64'h0E20000000000000;
    #10 assign a = 64'h2E9FFFFFFFFFFFFF; assign b = 64'h0E2FFFFFFFFFFFFF;

    #10 $display("\n2**-277 * 2**-798:");
    #10 assign a = 64'h2EA0000000000000; assign b = 64'h0E10000000000000;
    #10 assign a = 64'h2EAFFFFFFFFFFFFF; assign b = 64'h0E1FFFFFFFFFFFFF;

    #10 $display("\n2**-276 * 2**-799:");
    #10 assign a = 64'h2EB0000000000000; assign b = 64'h0E00000000000000;
    #10 assign a = 64'h2EBFFFFFFFFFFFFF; assign b = 64'h0E0FFFFFFFFFFFFF;

    #10 $display("\n2**-275 * 2**-800:");
    #10 assign a = 64'h2EC0000000000000; assign b = 64'h0DF0000000000000;
    #10 assign a = 64'h2ECFFFFFFFFFFFFF; assign b = 64'h0DFFFFFFFFFFFFFF;

    #10 $display("\n2**-274 * 2**-801:");
    #10 assign a = 64'h2ED0000000000000; assign b = 64'h0DE0000000000000;
    #10 assign a = 64'h2EDFFFFFFFFFFFFF; assign b = 64'h0DEFFFFFFFFFFFFF;

    #10 $display("\n2**-273 * 2**-802:");
    #10 assign a = 64'h2EE0000000000000; assign b = 64'h0DD0000000000000;
    #10 assign a = 64'h2EEFFFFFFFFFFFFF; assign b = 64'h0DDFFFFFFFFFFFFF;

    #10 $display("\n2**-272 * 2**-803:");
    #10 assign a = 64'h2EF0000000000000; assign b = 64'h0DC0000000000000;
    #10 assign a = 64'h2EFFFFFFFFFFFFFF; assign b = 64'h0DCFFFFFFFFFFFFF;

    #10 $display("\n2**-271 * 2**-804:");
    #10 assign a = 64'h2F00000000000000; assign b = 64'h0DB0000000000000;
    #10 assign a = 64'h2F0FFFFFFFFFFFFF; assign b = 64'h0DBFFFFFFFFFFFFF;

    #10 $display("\n2**-270 * 2**-805:");
    #10 assign a = 64'h2F10000000000000; assign b = 64'h0DA0000000000000;
    #10 assign a = 64'h2F1FFFFFFFFFFFFF; assign b = 64'h0DAFFFFFFFFFFFFF;

    #10 $display("\n2**-269 * 2**-806:");
    #10 assign a = 64'h2F20000000000000; assign b = 64'h0D90000000000000;
    #10 assign a = 64'h2F2FFFFFFFFFFFFF; assign b = 64'h0D9FFFFFFFFFFFFF;

    #10 $display("\n2**-268 * 2**-807:");
    #10 assign a = 64'h2F30000000000000; assign b = 64'h0D80000000000000;
    #10 assign a = 64'h2F3FFFFFFFFFFFFF; assign b = 64'h0D8FFFFFFFFFFFFF;

    #10 $display("\n2**-267 * 2**-808:");
    #10 assign a = 64'h2F40000000000000; assign b = 64'h0D70000000000000;
    #10 assign a = 64'h2F4FFFFFFFFFFFFF; assign b = 64'h0D7FFFFFFFFFFFFF;

    #10 $display("\n2**-266 * 2**-809:");
    #10 assign a = 64'h2F50000000000000; assign b = 64'h0D60000000000000;
    #10 assign a = 64'h2F5FFFFFFFFFFFFF; assign b = 64'h0D6FFFFFFFFFFFFF;

    #10 $display("\n2**-265 * 2**-810:");
    #10 assign a = 64'h2F60000000000000; assign b = 64'h0D50000000000000;
    #10 assign a = 64'h2F6FFFFFFFFFFFFF; assign b = 64'h0D5FFFFFFFFFFFFF;

    #10 $display("\n2**-264 * 2**-811:");
    #10 assign a = 64'h2F70000000000000; assign b = 64'h0D40000000000000;
    #10 assign a = 64'h2F7FFFFFFFFFFFFF; assign b = 64'h0D4FFFFFFFFFFFFF;

    #10 $display("\n2**-263 * 2**-812:");
    #10 assign a = 64'h2F80000000000000; assign b = 64'h0D30000000000000;
    #10 assign a = 64'h2F8FFFFFFFFFFFFF; assign b = 64'h0D3FFFFFFFFFFFFF;

    #10 $display("\n2**-262 * 2**-813:");
    #10 assign a = 64'h2F90000000000000; assign b = 64'h0D20000000000000;
    #10 assign a = 64'h2F9FFFFFFFFFFFFF; assign b = 64'h0D2FFFFFFFFFFFFF;

    #10 $display("\n2**-261 * 2**-814:");
    #10 assign a = 64'h2FA0000000000000; assign b = 64'h0D10000000000000;
    #10 assign a = 64'h2FAFFFFFFFFFFFFF; assign b = 64'h0D1FFFFFFFFFFFFF;

    #10 $display("\n2**-260 * 2**-815:");
    #10 assign a = 64'h2FB0000000000000; assign b = 64'h0D00000000000000;
    #10 assign a = 64'h2FBFFFFFFFFFFFFF; assign b = 64'h0D0FFFFFFFFFFFFF;

    #10 $display("\n2**-259 * 2**-816:");
    #10 assign a = 64'h2FC0000000000000; assign b = 64'h0CF0000000000000;
    #10 assign a = 64'h2FCFFFFFFFFFFFFF; assign b = 64'h0CFFFFFFFFFFFFFF;

    #10 $display("\n2**-258 * 2**-817:");
    #10 assign a = 64'h2FD0000000000000; assign b = 64'h0CE0000000000000;
    #10 assign a = 64'h2FDFFFFFFFFFFFFF; assign b = 64'h0CEFFFFFFFFFFFFF;

    #10 $display("\n2**-257 * 2**-818:");
    #10 assign a = 64'h2FE0000000000000; assign b = 64'h0CD0000000000000;
    #10 assign a = 64'h2FEFFFFFFFFFFFFF; assign b = 64'h0CDFFFFFFFFFFFFF;

    #10 $display("\n2**-256 * 2**-819:");
    #10 assign a = 64'h2FF0000000000000; assign b = 64'h0CC0000000000000;
    #10 assign a = 64'h2FFFFFFFFFFFFFFF; assign b = 64'h0CCFFFFFFFFFFFFF;

    #10 $display("\n2**-255 * 2**-820:");
    #10 assign a = 64'h3000000000000000; assign b = 64'h0CB0000000000000;
    #10 assign a = 64'h300FFFFFFFFFFFFF; assign b = 64'h0CBFFFFFFFFFFFFF;

    #10 $display("\n2**-254 * 2**-821:");
    #10 assign a = 64'h3010000000000000; assign b = 64'h0CA0000000000000;
    #10 assign a = 64'h301FFFFFFFFFFFFF; assign b = 64'h0CAFFFFFFFFFFFFF;

    #10 $display("\n2**-253 * 2**-822:");
    #10 assign a = 64'h3020000000000000; assign b = 64'h0C90000000000000;
    #10 assign a = 64'h302FFFFFFFFFFFFF; assign b = 64'h0C9FFFFFFFFFFFFF;

    #10 $display("\n2**-252 * 2**-823:");
    #10 assign a = 64'h3030000000000000; assign b = 64'h0C80000000000000;
    #10 assign a = 64'h303FFFFFFFFFFFFF; assign b = 64'h0C8FFFFFFFFFFFFF;

    #10 $display("\n2**-251 * 2**-824:");
    #10 assign a = 64'h3040000000000000; assign b = 64'h0C70000000000000;
    #10 assign a = 64'h304FFFFFFFFFFFFF; assign b = 64'h0C7FFFFFFFFFFFFF;

    #10 $display("\n2**-250 * 2**-825:");
    #10 assign a = 64'h3050000000000000; assign b = 64'h0C60000000000000;
    #10 assign a = 64'h305FFFFFFFFFFFFF; assign b = 64'h0C6FFFFFFFFFFFFF;

    #10 $display("\n2**-249 * 2**-826:");
    #10 assign a = 64'h3060000000000000; assign b = 64'h0C50000000000000;
    #10 assign a = 64'h306FFFFFFFFFFFFF; assign b = 64'h0C5FFFFFFFFFFFFF;

    #10 $display("\n2**-248 * 2**-827:");
    #10 assign a = 64'h3070000000000000; assign b = 64'h0C40000000000000;
    #10 assign a = 64'h307FFFFFFFFFFFFF; assign b = 64'h0C4FFFFFFFFFFFFF;

    #10 $display("\n2**-247 * 2**-828:");
    #10 assign a = 64'h3080000000000000; assign b = 64'h0C30000000000000;
    #10 assign a = 64'h308FFFFFFFFFFFFF; assign b = 64'h0C3FFFFFFFFFFFFF;

    #10 $display("\n2**-246 * 2**-829:");
    #10 assign a = 64'h3090000000000000; assign b = 64'h0C20000000000000;
    #10 assign a = 64'h309FFFFFFFFFFFFF; assign b = 64'h0C2FFFFFFFFFFFFF;

    #10 $display("\n2**-245 * 2**-830:");
    #10 assign a = 64'h30A0000000000000; assign b = 64'h0C10000000000000;
    #10 assign a = 64'h30AFFFFFFFFFFFFF; assign b = 64'h0C1FFFFFFFFFFFFF;

    #10 $display("\n2**-244 * 2**-831:");
    #10 assign a = 64'h30B0000000000000; assign b = 64'h0C00000000000000;
    #10 assign a = 64'h30BFFFFFFFFFFFFF; assign b = 64'h0C0FFFFFFFFFFFFF;

    #10 $display("\n2**-243 * 2**-832:");
    #10 assign a = 64'h30C0000000000000; assign b = 64'h0BF0000000000000;
    #10 assign a = 64'h30CFFFFFFFFFFFFF; assign b = 64'h0BFFFFFFFFFFFFFF;

    #10 $display("\n2**-242 * 2**-833:");
    #10 assign a = 64'h30D0000000000000; assign b = 64'h0BE0000000000000;
    #10 assign a = 64'h30DFFFFFFFFFFFFF; assign b = 64'h0BEFFFFFFFFFFFFF;

    #10 $display("\n2**-241 * 2**-834:");
    #10 assign a = 64'h30E0000000000000; assign b = 64'h0BD0000000000000;
    #10 assign a = 64'h30EFFFFFFFFFFFFF; assign b = 64'h0BDFFFFFFFFFFFFF;

    #10 $display("\n2**-240 * 2**-835:");
    #10 assign a = 64'h30F0000000000000; assign b = 64'h0BC0000000000000;
    #10 assign a = 64'h30FFFFFFFFFFFFFF; assign b = 64'h0BCFFFFFFFFFFFFF;

    #10 $display("\n2**-239 * 2**-836:");
    #10 assign a = 64'h3100000000000000; assign b = 64'h0BB0000000000000;
    #10 assign a = 64'h310FFFFFFFFFFFFF; assign b = 64'h0BBFFFFFFFFFFFFF;

    #10 $display("\n2**-238 * 2**-837:");
    #10 assign a = 64'h3110000000000000; assign b = 64'h0BA0000000000000;
    #10 assign a = 64'h311FFFFFFFFFFFFF; assign b = 64'h0BAFFFFFFFFFFFFF;

    #10 $display("\n2**-237 * 2**-838:");
    #10 assign a = 64'h3120000000000000; assign b = 64'h0B90000000000000;
    #10 assign a = 64'h312FFFFFFFFFFFFF; assign b = 64'h0B9FFFFFFFFFFFFF;

    #10 $display("\n2**-236 * 2**-839:");
    #10 assign a = 64'h3130000000000000; assign b = 64'h0B80000000000000;
    #10 assign a = 64'h313FFFFFFFFFFFFF; assign b = 64'h0B8FFFFFFFFFFFFF;

    #10 $display("\n2**-235 * 2**-840:");
    #10 assign a = 64'h3140000000000000; assign b = 64'h0B70000000000000;
    #10 assign a = 64'h314FFFFFFFFFFFFF; assign b = 64'h0B7FFFFFFFFFFFFF;

    #10 $display("\n2**-234 * 2**-841:");
    #10 assign a = 64'h3150000000000000; assign b = 64'h0B60000000000000;
    #10 assign a = 64'h315FFFFFFFFFFFFF; assign b = 64'h0B6FFFFFFFFFFFFF;

    #10 $display("\n2**-233 * 2**-842:");
    #10 assign a = 64'h3160000000000000; assign b = 64'h0B50000000000000;
    #10 assign a = 64'h316FFFFFFFFFFFFF; assign b = 64'h0B5FFFFFFFFFFFFF;

    #10 $display("\n2**-232 * 2**-843:");
    #10 assign a = 64'h3170000000000000; assign b = 64'h0B40000000000000;
    #10 assign a = 64'h317FFFFFFFFFFFFF; assign b = 64'h0B4FFFFFFFFFFFFF;

    #10 $display("\n2**-231 * 2**-844:");
    #10 assign a = 64'h3180000000000000; assign b = 64'h0B30000000000000;
    #10 assign a = 64'h318FFFFFFFFFFFFF; assign b = 64'h0B3FFFFFFFFFFFFF;

    #10 $display("\n2**-230 * 2**-845:");
    #10 assign a = 64'h3190000000000000; assign b = 64'h0B20000000000000;
    #10 assign a = 64'h319FFFFFFFFFFFFF; assign b = 64'h0B2FFFFFFFFFFFFF;

    #10 $display("\n2**-229 * 2**-846:");
    #10 assign a = 64'h31A0000000000000; assign b = 64'h0B10000000000000;
    #10 assign a = 64'h31AFFFFFFFFFFFFF; assign b = 64'h0B1FFFFFFFFFFFFF;

    #10 $display("\n2**-228 * 2**-847:");
    #10 assign a = 64'h31B0000000000000; assign b = 64'h0B00000000000000;
    #10 assign a = 64'h31BFFFFFFFFFFFFF; assign b = 64'h0B0FFFFFFFFFFFFF;

    #10 $display("\n2**-227 * 2**-848:");
    #10 assign a = 64'h31C0000000000000; assign b = 64'h0AF0000000000000;
    #10 assign a = 64'h31CFFFFFFFFFFFFF; assign b = 64'h0AFFFFFFFFFFFFFF;

    #10 $display("\n2**-226 * 2**-849:");
    #10 assign a = 64'h31D0000000000000; assign b = 64'h0AE0000000000000;
    #10 assign a = 64'h31DFFFFFFFFFFFFF; assign b = 64'h0AEFFFFFFFFFFFFF;

    #10 $display("\n2**-225 * 2**-850:");
    #10 assign a = 64'h31E0000000000000; assign b = 64'h0AD0000000000000;
    #10 assign a = 64'h31EFFFFFFFFFFFFF; assign b = 64'h0ADFFFFFFFFFFFFF;

    #10 $display("\n2**-224 * 2**-851:");
    #10 assign a = 64'h31F0000000000000; assign b = 64'h0AC0000000000000;
    #10 assign a = 64'h31FFFFFFFFFFFFFF; assign b = 64'h0ACFFFFFFFFFFFFF;

    #10 $display("\n2**-223 * 2**-852:");
    #10 assign a = 64'h3200000000000000; assign b = 64'h0AB0000000000000;
    #10 assign a = 64'h320FFFFFFFFFFFFF; assign b = 64'h0ABFFFFFFFFFFFFF;

    #10 $display("\n2**-222 * 2**-853:");
    #10 assign a = 64'h3210000000000000; assign b = 64'h0AA0000000000000;
    #10 assign a = 64'h321FFFFFFFFFFFFF; assign b = 64'h0AAFFFFFFFFFFFFF;

    #10 $display("\n2**-221 * 2**-854:");
    #10 assign a = 64'h3220000000000000; assign b = 64'h0A90000000000000;
    #10 assign a = 64'h322FFFFFFFFFFFFF; assign b = 64'h0A9FFFFFFFFFFFFF;

    #10 $display("\n2**-220 * 2**-855:");
    #10 assign a = 64'h3230000000000000; assign b = 64'h0A80000000000000;
    #10 assign a = 64'h323FFFFFFFFFFFFF; assign b = 64'h0A8FFFFFFFFFFFFF;

    #10 $display("\n2**-219 * 2**-856:");
    #10 assign a = 64'h3240000000000000; assign b = 64'h0A70000000000000;
    #10 assign a = 64'h324FFFFFFFFFFFFF; assign b = 64'h0A7FFFFFFFFFFFFF;

    #10 $display("\n2**-218 * 2**-857:");
    #10 assign a = 64'h3250000000000000; assign b = 64'h0A60000000000000;
    #10 assign a = 64'h325FFFFFFFFFFFFF; assign b = 64'h0A6FFFFFFFFFFFFF;

    #10 $display("\n2**-217 * 2**-858:");
    #10 assign a = 64'h3260000000000000; assign b = 64'h0A50000000000000;
    #10 assign a = 64'h326FFFFFFFFFFFFF; assign b = 64'h0A5FFFFFFFFFFFFF;

    #10 $display("\n2**-216 * 2**-859:");
    #10 assign a = 64'h3270000000000000; assign b = 64'h0A40000000000000;
    #10 assign a = 64'h327FFFFFFFFFFFFF; assign b = 64'h0A4FFFFFFFFFFFFF;

    #10 $display("\n2**-215 * 2**-860:");
    #10 assign a = 64'h3280000000000000; assign b = 64'h0A30000000000000;
    #10 assign a = 64'h328FFFFFFFFFFFFF; assign b = 64'h0A3FFFFFFFFFFFFF;

    #10 $display("\n2**-214 * 2**-861:");
    #10 assign a = 64'h3290000000000000; assign b = 64'h0A20000000000000;
    #10 assign a = 64'h329FFFFFFFFFFFFF; assign b = 64'h0A2FFFFFFFFFFFFF;

    #10 $display("\n2**-213 * 2**-862:");
    #10 assign a = 64'h32A0000000000000; assign b = 64'h0A10000000000000;
    #10 assign a = 64'h32AFFFFFFFFFFFFF; assign b = 64'h0A1FFFFFFFFFFFFF;

    #10 $display("\n2**-212 * 2**-863:");
    #10 assign a = 64'h32B0000000000000; assign b = 64'h0A00000000000000;
    #10 assign a = 64'h32BFFFFFFFFFFFFF; assign b = 64'h0A0FFFFFFFFFFFFF;

    #10 $display("\n2**-211 * 2**-864:");
    #10 assign a = 64'h32C0000000000000; assign b = 64'h09F0000000000000;
    #10 assign a = 64'h32CFFFFFFFFFFFFF; assign b = 64'h09FFFFFFFFFFFFFF;

    #10 $display("\n2**-210 * 2**-865:");
    #10 assign a = 64'h32D0000000000000; assign b = 64'h09E0000000000000;
    #10 assign a = 64'h32DFFFFFFFFFFFFF; assign b = 64'h09EFFFFFFFFFFFFF;

    #10 $display("\n2**-209 * 2**-866:");
    #10 assign a = 64'h32E0000000000000; assign b = 64'h09D0000000000000;
    #10 assign a = 64'h32EFFFFFFFFFFFFF; assign b = 64'h09DFFFFFFFFFFFFF;

    #10 $display("\n2**-208 * 2**-867:");
    #10 assign a = 64'h32F0000000000000; assign b = 64'h09C0000000000000;
    #10 assign a = 64'h32FFFFFFFFFFFFFF; assign b = 64'h09CFFFFFFFFFFFFF;

    #10 $display("\n2**-207 * 2**-868:");
    #10 assign a = 64'h3300000000000000; assign b = 64'h09B0000000000000;
    #10 assign a = 64'h330FFFFFFFFFFFFF; assign b = 64'h09BFFFFFFFFFFFFF;

    #10 $display("\n2**-206 * 2**-869:");
    #10 assign a = 64'h3310000000000000; assign b = 64'h09A0000000000000;
    #10 assign a = 64'h331FFFFFFFFFFFFF; assign b = 64'h09AFFFFFFFFFFFFF;

    #10 $display("\n2**-205 * 2**-870:");
    #10 assign a = 64'h3320000000000000; assign b = 64'h0990000000000000;
    #10 assign a = 64'h332FFFFFFFFFFFFF; assign b = 64'h099FFFFFFFFFFFFF;

    #10 $display("\n2**-204 * 2**-871:");
    #10 assign a = 64'h3330000000000000; assign b = 64'h0980000000000000;
    #10 assign a = 64'h333FFFFFFFFFFFFF; assign b = 64'h098FFFFFFFFFFFFF;

    #10 $display("\n2**-203 * 2**-872:");
    #10 assign a = 64'h3340000000000000; assign b = 64'h0970000000000000;
    #10 assign a = 64'h334FFFFFFFFFFFFF; assign b = 64'h097FFFFFFFFFFFFF;

    #10 $display("\n2**-202 * 2**-873:");
    #10 assign a = 64'h3350000000000000; assign b = 64'h0960000000000000;
    #10 assign a = 64'h335FFFFFFFFFFFFF; assign b = 64'h096FFFFFFFFFFFFF;

    #10 $display("\n2**-201 * 2**-874:");
    #10 assign a = 64'h3360000000000000; assign b = 64'h0950000000000000;
    #10 assign a = 64'h336FFFFFFFFFFFFF; assign b = 64'h095FFFFFFFFFFFFF;

    #10 $display("\n2**-200 * 2**-875:");
    #10 assign a = 64'h3370000000000000; assign b = 64'h0940000000000000;
    #10 assign a = 64'h337FFFFFFFFFFFFF; assign b = 64'h094FFFFFFFFFFFFF;

    #10 $display("\n2**-199 * 2**-876:");
    #10 assign a = 64'h3380000000000000; assign b = 64'h0930000000000000;
    #10 assign a = 64'h338FFFFFFFFFFFFF; assign b = 64'h093FFFFFFFFFFFFF;

    #10 $display("\n2**-198 * 2**-877:");
    #10 assign a = 64'h3390000000000000; assign b = 64'h0920000000000000;
    #10 assign a = 64'h339FFFFFFFFFFFFF; assign b = 64'h092FFFFFFFFFFFFF;

    #10 $display("\n2**-197 * 2**-878:");
    #10 assign a = 64'h33A0000000000000; assign b = 64'h0910000000000000;
    #10 assign a = 64'h33AFFFFFFFFFFFFF; assign b = 64'h091FFFFFFFFFFFFF;

    #10 $display("\n2**-196 * 2**-879:");
    #10 assign a = 64'h33B0000000000000; assign b = 64'h0900000000000000;
    #10 assign a = 64'h33BFFFFFFFFFFFFF; assign b = 64'h090FFFFFFFFFFFFF;

    #10 $display("\n2**-195 * 2**-880:");
    #10 assign a = 64'h33C0000000000000; assign b = 64'h08F0000000000000;
    #10 assign a = 64'h33CFFFFFFFFFFFFF; assign b = 64'h08FFFFFFFFFFFFFF;

    #10 $display("\n2**-194 * 2**-881:");
    #10 assign a = 64'h33D0000000000000; assign b = 64'h08E0000000000000;
    #10 assign a = 64'h33DFFFFFFFFFFFFF; assign b = 64'h08EFFFFFFFFFFFFF;

    #10 $display("\n2**-193 * 2**-882:");
    #10 assign a = 64'h33E0000000000000; assign b = 64'h08D0000000000000;
    #10 assign a = 64'h33EFFFFFFFFFFFFF; assign b = 64'h08DFFFFFFFFFFFFF;

    #10 $display("\n2**-192 * 2**-883:");
    #10 assign a = 64'h33F0000000000000; assign b = 64'h08C0000000000000;
    #10 assign a = 64'h33FFFFFFFFFFFFFF; assign b = 64'h08CFFFFFFFFFFFFF;

    #10 $display("\n2**-191 * 2**-884:");
    #10 assign a = 64'h3400000000000000; assign b = 64'h08B0000000000000;
    #10 assign a = 64'h340FFFFFFFFFFFFF; assign b = 64'h08BFFFFFFFFFFFFF;

    #10 $display("\n2**-190 * 2**-885:");
    #10 assign a = 64'h3410000000000000; assign b = 64'h08A0000000000000;
    #10 assign a = 64'h341FFFFFFFFFFFFF; assign b = 64'h08AFFFFFFFFFFFFF;

    #10 $display("\n2**-189 * 2**-886:");
    #10 assign a = 64'h3420000000000000; assign b = 64'h0890000000000000;
    #10 assign a = 64'h342FFFFFFFFFFFFF; assign b = 64'h089FFFFFFFFFFFFF;

    #10 $display("\n2**-188 * 2**-887:");
    #10 assign a = 64'h3430000000000000; assign b = 64'h0880000000000000;
    #10 assign a = 64'h343FFFFFFFFFFFFF; assign b = 64'h088FFFFFFFFFFFFF;

    #10 $display("\n2**-187 * 2**-888:");
    #10 assign a = 64'h3440000000000000; assign b = 64'h0870000000000000;
    #10 assign a = 64'h344FFFFFFFFFFFFF; assign b = 64'h087FFFFFFFFFFFFF;

    #10 $display("\n2**-186 * 2**-889:");
    #10 assign a = 64'h3450000000000000; assign b = 64'h0860000000000000;
    #10 assign a = 64'h345FFFFFFFFFFFFF; assign b = 64'h086FFFFFFFFFFFFF;

    #10 $display("\n2**-185 * 2**-890:");
    #10 assign a = 64'h3460000000000000; assign b = 64'h0850000000000000;
    #10 assign a = 64'h346FFFFFFFFFFFFF; assign b = 64'h085FFFFFFFFFFFFF;

    #10 $display("\n2**-184 * 2**-891:");
    #10 assign a = 64'h3470000000000000; assign b = 64'h0840000000000000;
    #10 assign a = 64'h347FFFFFFFFFFFFF; assign b = 64'h084FFFFFFFFFFFFF;

    #10 $display("\n2**-183 * 2**-892:");
    #10 assign a = 64'h3480000000000000; assign b = 64'h0830000000000000;
    #10 assign a = 64'h348FFFFFFFFFFFFF; assign b = 64'h083FFFFFFFFFFFFF;

    #10 $display("\n2**-182 * 2**-893:");
    #10 assign a = 64'h3490000000000000; assign b = 64'h0820000000000000;
    #10 assign a = 64'h349FFFFFFFFFFFFF; assign b = 64'h082FFFFFFFFFFFFF;

    #10 $display("\n2**-181 * 2**-894:");
    #10 assign a = 64'h34A0000000000000; assign b = 64'h0810000000000000;
    #10 assign a = 64'h34AFFFFFFFFFFFFF; assign b = 64'h081FFFFFFFFFFFFF;

    #10 $display("\n2**-180 * 2**-895:");
    #10 assign a = 64'h34B0000000000000; assign b = 64'h0800000000000000;
    #10 assign a = 64'h34BFFFFFFFFFFFFF; assign b = 64'h080FFFFFFFFFFFFF;

    #10 $display("\n2**-179 * 2**-896:");
    #10 assign a = 64'h34C0000000000000; assign b = 64'h07F0000000000000;
    #10 assign a = 64'h34CFFFFFFFFFFFFF; assign b = 64'h07FFFFFFFFFFFFFF;

    #10 $display("\n2**-178 * 2**-897:");
    #10 assign a = 64'h34D0000000000000; assign b = 64'h07E0000000000000;
    #10 assign a = 64'h34DFFFFFFFFFFFFF; assign b = 64'h07EFFFFFFFFFFFFF;

    #10 $display("\n2**-177 * 2**-898:");
    #10 assign a = 64'h34E0000000000000; assign b = 64'h07D0000000000000;
    #10 assign a = 64'h34EFFFFFFFFFFFFF; assign b = 64'h07DFFFFFFFFFFFFF;

    #10 $display("\n2**-176 * 2**-899:");
    #10 assign a = 64'h34F0000000000000; assign b = 64'h07C0000000000000;
    #10 assign a = 64'h34FFFFFFFFFFFFFF; assign b = 64'h07CFFFFFFFFFFFFF;

    #10 $display("\n2**-175 * 2**-900:");
    #10 assign a = 64'h3500000000000000; assign b = 64'h07B0000000000000;
    #10 assign a = 64'h350FFFFFFFFFFFFF; assign b = 64'h07BFFFFFFFFFFFFF;

    #10 $display("\n2**-174 * 2**-901:");
    #10 assign a = 64'h3510000000000000; assign b = 64'h07A0000000000000;
    #10 assign a = 64'h351FFFFFFFFFFFFF; assign b = 64'h07AFFFFFFFFFFFFF;

    #10 $display("\n2**-173 * 2**-902:");
    #10 assign a = 64'h3520000000000000; assign b = 64'h0790000000000000;
    #10 assign a = 64'h352FFFFFFFFFFFFF; assign b = 64'h079FFFFFFFFFFFFF;

    #10 $display("\n2**-172 * 2**-903:");
    #10 assign a = 64'h3530000000000000; assign b = 64'h0780000000000000;
    #10 assign a = 64'h353FFFFFFFFFFFFF; assign b = 64'h078FFFFFFFFFFFFF;

    #10 $display("\n2**-171 * 2**-904:");
    #10 assign a = 64'h3540000000000000; assign b = 64'h0770000000000000;
    #10 assign a = 64'h354FFFFFFFFFFFFF; assign b = 64'h077FFFFFFFFFFFFF;

    #10 $display("\n2**-170 * 2**-905:");
    #10 assign a = 64'h3550000000000000; assign b = 64'h0760000000000000;
    #10 assign a = 64'h355FFFFFFFFFFFFF; assign b = 64'h076FFFFFFFFFFFFF;

    #10 $display("\n2**-169 * 2**-906:");
    #10 assign a = 64'h3560000000000000; assign b = 64'h0750000000000000;
    #10 assign a = 64'h356FFFFFFFFFFFFF; assign b = 64'h075FFFFFFFFFFFFF;

    #10 $display("\n2**-168 * 2**-907:");
    #10 assign a = 64'h3570000000000000; assign b = 64'h0740000000000000;
    #10 assign a = 64'h357FFFFFFFFFFFFF; assign b = 64'h074FFFFFFFFFFFFF;

    #10 $display("\n2**-167 * 2**-908:");
    #10 assign a = 64'h3580000000000000; assign b = 64'h0730000000000000;
    #10 assign a = 64'h358FFFFFFFFFFFFF; assign b = 64'h073FFFFFFFFFFFFF;

    #10 $display("\n2**-166 * 2**-909:");
    #10 assign a = 64'h3590000000000000; assign b = 64'h0720000000000000;
    #10 assign a = 64'h359FFFFFFFFFFFFF; assign b = 64'h072FFFFFFFFFFFFF;

    #10 $display("\n2**-165 * 2**-910:");
    #10 assign a = 64'h35A0000000000000; assign b = 64'h0710000000000000;
    #10 assign a = 64'h35AFFFFFFFFFFFFF; assign b = 64'h071FFFFFFFFFFFFF;

    #10 $display("\n2**-164 * 2**-911:");
    #10 assign a = 64'h35B0000000000000; assign b = 64'h0700000000000000;
    #10 assign a = 64'h35BFFFFFFFFFFFFF; assign b = 64'h070FFFFFFFFFFFFF;

    #10 $display("\n2**-163 * 2**-912:");
    #10 assign a = 64'h35C0000000000000; assign b = 64'h06F0000000000000;
    #10 assign a = 64'h35CFFFFFFFFFFFFF; assign b = 64'h06FFFFFFFFFFFFFF;

    #10 $display("\n2**-162 * 2**-913:");
    #10 assign a = 64'h35D0000000000000; assign b = 64'h06E0000000000000;
    #10 assign a = 64'h35DFFFFFFFFFFFFF; assign b = 64'h06EFFFFFFFFFFFFF;

    #10 $display("\n2**-161 * 2**-914:");
    #10 assign a = 64'h35E0000000000000; assign b = 64'h06D0000000000000;
    #10 assign a = 64'h35EFFFFFFFFFFFFF; assign b = 64'h06DFFFFFFFFFFFFF;

    #10 $display("\n2**-160 * 2**-915:");
    #10 assign a = 64'h35F0000000000000; assign b = 64'h06C0000000000000;
    #10 assign a = 64'h35FFFFFFFFFFFFFF; assign b = 64'h06CFFFFFFFFFFFFF;

    #10 $display("\n2**-159 * 2**-916:");
    #10 assign a = 64'h3600000000000000; assign b = 64'h06B0000000000000;
    #10 assign a = 64'h360FFFFFFFFFFFFF; assign b = 64'h06BFFFFFFFFFFFFF;

    #10 $display("\n2**-158 * 2**-917:");
    #10 assign a = 64'h3610000000000000; assign b = 64'h06A0000000000000;
    #10 assign a = 64'h361FFFFFFFFFFFFF; assign b = 64'h06AFFFFFFFFFFFFF;

    #10 $display("\n2**-157 * 2**-918:");
    #10 assign a = 64'h3620000000000000; assign b = 64'h0690000000000000;
    #10 assign a = 64'h362FFFFFFFFFFFFF; assign b = 64'h069FFFFFFFFFFFFF;

    #10 $display("\n2**-156 * 2**-919:");
    #10 assign a = 64'h3630000000000000; assign b = 64'h0680000000000000;
    #10 assign a = 64'h363FFFFFFFFFFFFF; assign b = 64'h068FFFFFFFFFFFFF;

    #10 $display("\n2**-155 * 2**-920:");
    #10 assign a = 64'h3640000000000000; assign b = 64'h0670000000000000;
    #10 assign a = 64'h364FFFFFFFFFFFFF; assign b = 64'h067FFFFFFFFFFFFF;

    #10 $display("\n2**-154 * 2**-921:");
    #10 assign a = 64'h3650000000000000; assign b = 64'h0660000000000000;
    #10 assign a = 64'h365FFFFFFFFFFFFF; assign b = 64'h066FFFFFFFFFFFFF;

    #10 $display("\n2**-153 * 2**-922:");
    #10 assign a = 64'h3660000000000000; assign b = 64'h0650000000000000;
    #10 assign a = 64'h366FFFFFFFFFFFFF; assign b = 64'h065FFFFFFFFFFFFF;

    #10 $display("\n2**-152 * 2**-923:");
    #10 assign a = 64'h3670000000000000; assign b = 64'h0640000000000000;
    #10 assign a = 64'h367FFFFFFFFFFFFF; assign b = 64'h064FFFFFFFFFFFFF;

    #10 $display("\n2**-151 * 2**-924:");
    #10 assign a = 64'h3680000000000000; assign b = 64'h0630000000000000;
    #10 assign a = 64'h368FFFFFFFFFFFFF; assign b = 64'h063FFFFFFFFFFFFF;

    #10 $display("\n2**-150 * 2**-925:");
    #10 assign a = 64'h3690000000000000; assign b = 64'h0620000000000000;
    #10 assign a = 64'h369FFFFFFFFFFFFF; assign b = 64'h062FFFFFFFFFFFFF;

    #10 $display("\n2**-149 * 2**-926:");
    #10 assign a = 64'h36A0000000000000; assign b = 64'h0610000000000000;
    #10 assign a = 64'h36AFFFFFFFFFFFFF; assign b = 64'h061FFFFFFFFFFFFF;

    #10 $display("\n2**-148 * 2**-927:");
    #10 assign a = 64'h36B0000000000000; assign b = 64'h0600000000000000;
    #10 assign a = 64'h36BFFFFFFFFFFFFF; assign b = 64'h060FFFFFFFFFFFFF;

    #10 $display("\n2**-147 * 2**-928:");
    #10 assign a = 64'h36C0000000000000; assign b = 64'h05F0000000000000;
    #10 assign a = 64'h36CFFFFFFFFFFFFF; assign b = 64'h05FFFFFFFFFFFFFF;

    #10 $display("\n2**-146 * 2**-929:");
    #10 assign a = 64'h36D0000000000000; assign b = 64'h05E0000000000000;
    #10 assign a = 64'h36DFFFFFFFFFFFFF; assign b = 64'h05EFFFFFFFFFFFFF;

    #10 $display("\n2**-145 * 2**-930:");
    #10 assign a = 64'h36E0000000000000; assign b = 64'h05D0000000000000;
    #10 assign a = 64'h36EFFFFFFFFFFFFF; assign b = 64'h05DFFFFFFFFFFFFF;

    #10 $display("\n2**-144 * 2**-931:");
    #10 assign a = 64'h36F0000000000000; assign b = 64'h05C0000000000000;
    #10 assign a = 64'h36FFFFFFFFFFFFFF; assign b = 64'h05CFFFFFFFFFFFFF;

    #10 $display("\n2**-143 * 2**-932:");
    #10 assign a = 64'h3700000000000000; assign b = 64'h05B0000000000000;
    #10 assign a = 64'h370FFFFFFFFFFFFF; assign b = 64'h05BFFFFFFFFFFFFF;

    #10 $display("\n2**-142 * 2**-933:");
    #10 assign a = 64'h3710000000000000; assign b = 64'h05A0000000000000;
    #10 assign a = 64'h371FFFFFFFFFFFFF; assign b = 64'h05AFFFFFFFFFFFFF;

    #10 $display("\n2**-141 * 2**-934:");
    #10 assign a = 64'h3720000000000000; assign b = 64'h0590000000000000;
    #10 assign a = 64'h372FFFFFFFFFFFFF; assign b = 64'h059FFFFFFFFFFFFF;

    #10 $display("\n2**-140 * 2**-935:");
    #10 assign a = 64'h3730000000000000; assign b = 64'h0580000000000000;
    #10 assign a = 64'h373FFFFFFFFFFFFF; assign b = 64'h058FFFFFFFFFFFFF;

    #10 $display("\n2**-139 * 2**-936:");
    #10 assign a = 64'h3740000000000000; assign b = 64'h0570000000000000;
    #10 assign a = 64'h374FFFFFFFFFFFFF; assign b = 64'h057FFFFFFFFFFFFF;

    #10 $display("\n2**-138 * 2**-937:");
    #10 assign a = 64'h3750000000000000; assign b = 64'h0560000000000000;
    #10 assign a = 64'h375FFFFFFFFFFFFF; assign b = 64'h056FFFFFFFFFFFFF;

    #10 $display("\n2**-137 * 2**-938:");
    #10 assign a = 64'h3760000000000000; assign b = 64'h0550000000000000;
    #10 assign a = 64'h376FFFFFFFFFFFFF; assign b = 64'h055FFFFFFFFFFFFF;

    #10 $display("\n2**-136 * 2**-939:");
    #10 assign a = 64'h3770000000000000; assign b = 64'h0540000000000000;
    #10 assign a = 64'h377FFFFFFFFFFFFF; assign b = 64'h054FFFFFFFFFFFFF;

    #10 $display("\n2**-135 * 2**-940:");
    #10 assign a = 64'h3780000000000000; assign b = 64'h0530000000000000;
    #10 assign a = 64'h378FFFFFFFFFFFFF; assign b = 64'h053FFFFFFFFFFFFF;

    #10 $display("\n2**-134 * 2**-941:");
    #10 assign a = 64'h3790000000000000; assign b = 64'h0520000000000000;
    #10 assign a = 64'h379FFFFFFFFFFFFF; assign b = 64'h052FFFFFFFFFFFFF;

    #10 $display("\n2**-133 * 2**-942:");
    #10 assign a = 64'h37A0000000000000; assign b = 64'h0510000000000000;
    #10 assign a = 64'h37AFFFFFFFFFFFFF; assign b = 64'h051FFFFFFFFFFFFF;

    #10 $display("\n2**-132 * 2**-943:");
    #10 assign a = 64'h37B0000000000000; assign b = 64'h0500000000000000;
    #10 assign a = 64'h37BFFFFFFFFFFFFF; assign b = 64'h050FFFFFFFFFFFFF;

    #10 $display("\n2**-131 * 2**-944:");
    #10 assign a = 64'h37C0000000000000; assign b = 64'h04F0000000000000;
    #10 assign a = 64'h37CFFFFFFFFFFFFF; assign b = 64'h04FFFFFFFFFFFFFF;

    #10 $display("\n2**-130 * 2**-945:");
    #10 assign a = 64'h37D0000000000000; assign b = 64'h04E0000000000000;
    #10 assign a = 64'h37DFFFFFFFFFFFFF; assign b = 64'h04EFFFFFFFFFFFFF;

    #10 $display("\n2**-129 * 2**-946:");
    #10 assign a = 64'h37E0000000000000; assign b = 64'h04D0000000000000;
    #10 assign a = 64'h37EFFFFFFFFFFFFF; assign b = 64'h04DFFFFFFFFFFFFF;

    #10 $display("\n2**-128 * 2**-947:");
    #10 assign a = 64'h37F0000000000000; assign b = 64'h04C0000000000000;
    #10 assign a = 64'h37FFFFFFFFFFFFFF; assign b = 64'h04CFFFFFFFFFFFFF;

    #10 $display("\n2**-127 * 2**-948:");
    #10 assign a = 64'h3800000000000000; assign b = 64'h04B0000000000000;
    #10 assign a = 64'h380FFFFFFFFFFFFF; assign b = 64'h04BFFFFFFFFFFFFF;

    #10 $display("\n2**-126 * 2**-949:");
    #10 assign a = 64'h3810000000000000; assign b = 64'h04A0000000000000;
    #10 assign a = 64'h381FFFFFFFFFFFFF; assign b = 64'h04AFFFFFFFFFFFFF;

    #10 $display("\n2**-125 * 2**-950:");
    #10 assign a = 64'h3820000000000000; assign b = 64'h0490000000000000;
    #10 assign a = 64'h382FFFFFFFFFFFFF; assign b = 64'h049FFFFFFFFFFFFF;

    #10 $display("\n2**-124 * 2**-951:");
    #10 assign a = 64'h3830000000000000; assign b = 64'h0480000000000000;
    #10 assign a = 64'h383FFFFFFFFFFFFF; assign b = 64'h048FFFFFFFFFFFFF;

    #10 $display("\n2**-123 * 2**-952:");
    #10 assign a = 64'h3840000000000000; assign b = 64'h0470000000000000;
    #10 assign a = 64'h384FFFFFFFFFFFFF; assign b = 64'h047FFFFFFFFFFFFF;

    #10 $display("\n2**-122 * 2**-953:");
    #10 assign a = 64'h3850000000000000; assign b = 64'h0460000000000000;
    #10 assign a = 64'h385FFFFFFFFFFFFF; assign b = 64'h046FFFFFFFFFFFFF;

    #10 $display("\n2**-121 * 2**-954:");
    #10 assign a = 64'h3860000000000000; assign b = 64'h0450000000000000;
    #10 assign a = 64'h386FFFFFFFFFFFFF; assign b = 64'h045FFFFFFFFFFFFF;

    #10 $display("\n2**-120 * 2**-955:");
    #10 assign a = 64'h3870000000000000; assign b = 64'h0440000000000000;
    #10 assign a = 64'h387FFFFFFFFFFFFF; assign b = 64'h044FFFFFFFFFFFFF;

    #10 $display("\n2**-119 * 2**-956:");
    #10 assign a = 64'h3880000000000000; assign b = 64'h0430000000000000;
    #10 assign a = 64'h388FFFFFFFFFFFFF; assign b = 64'h043FFFFFFFFFFFFF;

    #10 $display("\n2**-118 * 2**-957:");
    #10 assign a = 64'h3890000000000000; assign b = 64'h0420000000000000;
    #10 assign a = 64'h389FFFFFFFFFFFFF; assign b = 64'h042FFFFFFFFFFFFF;

    #10 $display("\n2**-117 * 2**-958:");
    #10 assign a = 64'h38A0000000000000; assign b = 64'h0410000000000000;
    #10 assign a = 64'h38AFFFFFFFFFFFFF; assign b = 64'h041FFFFFFFFFFFFF;

    #10 $display("\n2**-116 * 2**-959:");
    #10 assign a = 64'h38B0000000000000; assign b = 64'h0400000000000000;
    #10 assign a = 64'h38BFFFFFFFFFFFFF; assign b = 64'h040FFFFFFFFFFFFF;

    #10 $display("\n2**-115 * 2**-960:");
    #10 assign a = 64'h38C0000000000000; assign b = 64'h03F0000000000000;
    #10 assign a = 64'h38CFFFFFFFFFFFFF; assign b = 64'h03FFFFFFFFFFFFFF;

    #10 $display("\n2**-114 * 2**-961:");
    #10 assign a = 64'h38D0000000000000; assign b = 64'h03E0000000000000;
    #10 assign a = 64'h38DFFFFFFFFFFFFF; assign b = 64'h03EFFFFFFFFFFFFF;

    #10 $display("\n2**-113 * 2**-962:");
    #10 assign a = 64'h38E0000000000000; assign b = 64'h03D0000000000000;
    #10 assign a = 64'h38EFFFFFFFFFFFFF; assign b = 64'h03DFFFFFFFFFFFFF;

    #10 $display("\n2**-112 * 2**-963:");
    #10 assign a = 64'h38F0000000000000; assign b = 64'h03C0000000000000;
    #10 assign a = 64'h38FFFFFFFFFFFFFF; assign b = 64'h03CFFFFFFFFFFFFF;

    #10 $display("\n2**-111 * 2**-964:");
    #10 assign a = 64'h3900000000000000; assign b = 64'h03B0000000000000;
    #10 assign a = 64'h390FFFFFFFFFFFFF; assign b = 64'h03BFFFFFFFFFFFFF;

    #10 $display("\n2**-110 * 2**-965:");
    #10 assign a = 64'h3910000000000000; assign b = 64'h03A0000000000000;
    #10 assign a = 64'h391FFFFFFFFFFFFF; assign b = 64'h03AFFFFFFFFFFFFF;

    #10 $display("\n2**-109 * 2**-966:");
    #10 assign a = 64'h3920000000000000; assign b = 64'h0390000000000000;
    #10 assign a = 64'h392FFFFFFFFFFFFF; assign b = 64'h039FFFFFFFFFFFFF;

    #10 $display("\n2**-108 * 2**-967:");
    #10 assign a = 64'h3930000000000000; assign b = 64'h0380000000000000;
    #10 assign a = 64'h393FFFFFFFFFFFFF; assign b = 64'h038FFFFFFFFFFFFF;

    #10 $display("\n2**-107 * 2**-968:");
    #10 assign a = 64'h3940000000000000; assign b = 64'h0370000000000000;
    #10 assign a = 64'h394FFFFFFFFFFFFF; assign b = 64'h037FFFFFFFFFFFFF;

    #10 $display("\n2**-106 * 2**-969:");
    #10 assign a = 64'h3950000000000000; assign b = 64'h0360000000000000;
    #10 assign a = 64'h395FFFFFFFFFFFFF; assign b = 64'h036FFFFFFFFFFFFF;

    #10 $display("\n2**-105 * 2**-970:");
    #10 assign a = 64'h3960000000000000; assign b = 64'h0350000000000000;
    #10 assign a = 64'h396FFFFFFFFFFFFF; assign b = 64'h035FFFFFFFFFFFFF;

    #10 $display("\n2**-104 * 2**-971:");
    #10 assign a = 64'h3970000000000000; assign b = 64'h0340000000000000;
    #10 assign a = 64'h397FFFFFFFFFFFFF; assign b = 64'h034FFFFFFFFFFFFF;

    #10 $display("\n2**-103 * 2**-972:");
    #10 assign a = 64'h3980000000000000; assign b = 64'h0330000000000000;
    #10 assign a = 64'h398FFFFFFFFFFFFF; assign b = 64'h033FFFFFFFFFFFFF;

    #10 $display("\n2**-102 * 2**-973:");
    #10 assign a = 64'h3990000000000000; assign b = 64'h0320000000000000;
    #10 assign a = 64'h399FFFFFFFFFFFFF; assign b = 64'h032FFFFFFFFFFFFF;

    #10 $display("\n2**-101 * 2**-974:");
    #10 assign a = 64'h39A0000000000000; assign b = 64'h0310000000000000;
    #10 assign a = 64'h39AFFFFFFFFFFFFF; assign b = 64'h031FFFFFFFFFFFFF;

    #10 $display("\n2**-100 * 2**-975:");
    #10 assign a = 64'h39B0000000000000; assign b = 64'h0300000000000000;
    #10 assign a = 64'h39BFFFFFFFFFFFFF; assign b = 64'h030FFFFFFFFFFFFF;

    #10 $display("\n2**-99 * 2**-976:");
    #10 assign a = 64'h39C0000000000000; assign b = 64'h02F0000000000000;
    #10 assign a = 64'h39CFFFFFFFFFFFFF; assign b = 64'h02FFFFFFFFFFFFFF;

    #10 $display("\n2**-98 * 2**-977:");
    #10 assign a = 64'h39D0000000000000; assign b = 64'h02E0000000000000;
    #10 assign a = 64'h39DFFFFFFFFFFFFF; assign b = 64'h02EFFFFFFFFFFFFF;

    #10 $display("\n2**-97 * 2**-978:");
    #10 assign a = 64'h39E0000000000000; assign b = 64'h02D0000000000000;
    #10 assign a = 64'h39EFFFFFFFFFFFFF; assign b = 64'h02DFFFFFFFFFFFFF;

    #10 $display("\n2**-96 * 2**-979:");
    #10 assign a = 64'h39F0000000000000; assign b = 64'h02C0000000000000;
    #10 assign a = 64'h39FFFFFFFFFFFFFF; assign b = 64'h02CFFFFFFFFFFFFF;

    #10 $display("\n2**-95 * 2**-980:");
    #10 assign a = 64'h3A00000000000000; assign b = 64'h02B0000000000000;
    #10 assign a = 64'h3A0FFFFFFFFFFFFF; assign b = 64'h02BFFFFFFFFFFFFF;

    #10 $display("\n2**-94 * 2**-981:");
    #10 assign a = 64'h3A10000000000000; assign b = 64'h02A0000000000000;
    #10 assign a = 64'h3A1FFFFFFFFFFFFF; assign b = 64'h02AFFFFFFFFFFFFF;

    #10 $display("\n2**-93 * 2**-982:");
    #10 assign a = 64'h3A20000000000000; assign b = 64'h0290000000000000;
    #10 assign a = 64'h3A2FFFFFFFFFFFFF; assign b = 64'h029FFFFFFFFFFFFF;

    #10 $display("\n2**-92 * 2**-983:");
    #10 assign a = 64'h3A30000000000000; assign b = 64'h0280000000000000;
    #10 assign a = 64'h3A3FFFFFFFFFFFFF; assign b = 64'h028FFFFFFFFFFFFF;

    #10 $display("\n2**-91 * 2**-984:");
    #10 assign a = 64'h3A40000000000000; assign b = 64'h0270000000000000;
    #10 assign a = 64'h3A4FFFFFFFFFFFFF; assign b = 64'h027FFFFFFFFFFFFF;

    #10 $display("\n2**-90 * 2**-985:");
    #10 assign a = 64'h3A50000000000000; assign b = 64'h0260000000000000;
    #10 assign a = 64'h3A5FFFFFFFFFFFFF; assign b = 64'h026FFFFFFFFFFFFF;

    #10 $display("\n2**-89 * 2**-986:");
    #10 assign a = 64'h3A60000000000000; assign b = 64'h0250000000000000;
    #10 assign a = 64'h3A6FFFFFFFFFFFFF; assign b = 64'h025FFFFFFFFFFFFF;

    #10 $display("\n2**-88 * 2**-987:");
    #10 assign a = 64'h3A70000000000000; assign b = 64'h0240000000000000;
    #10 assign a = 64'h3A7FFFFFFFFFFFFF; assign b = 64'h024FFFFFFFFFFFFF;

    #10 $display("\n2**-87 * 2**-988:");
    #10 assign a = 64'h3A80000000000000; assign b = 64'h0230000000000000;
    #10 assign a = 64'h3A8FFFFFFFFFFFFF; assign b = 64'h023FFFFFFFFFFFFF;

    #10 $display("\n2**-86 * 2**-989:");
    #10 assign a = 64'h3A90000000000000; assign b = 64'h0220000000000000;
    #10 assign a = 64'h3A9FFFFFFFFFFFFF; assign b = 64'h022FFFFFFFFFFFFF;

    #10 $display("\n2**-85 * 2**-990:");
    #10 assign a = 64'h3AA0000000000000; assign b = 64'h0210000000000000;
    #10 assign a = 64'h3AAFFFFFFFFFFFFF; assign b = 64'h021FFFFFFFFFFFFF;

    #10 $display("\n2**-84 * 2**-991:");
    #10 assign a = 64'h3AB0000000000000; assign b = 64'h0200000000000000;
    #10 assign a = 64'h3ABFFFFFFFFFFFFF; assign b = 64'h020FFFFFFFFFFFFF;

    #10 $display("\n2**-83 * 2**-992:");
    #10 assign a = 64'h3AC0000000000000; assign b = 64'h01F0000000000000;
    #10 assign a = 64'h3ACFFFFFFFFFFFFF; assign b = 64'h01FFFFFFFFFFFFFF;

    #10 $display("\n2**-82 * 2**-993:");
    #10 assign a = 64'h3AD0000000000000; assign b = 64'h01E0000000000000;
    #10 assign a = 64'h3ADFFFFFFFFFFFFF; assign b = 64'h01EFFFFFFFFFFFFF;

    #10 $display("\n2**-81 * 2**-994:");
    #10 assign a = 64'h3AE0000000000000; assign b = 64'h01D0000000000000;
    #10 assign a = 64'h3AEFFFFFFFFFFFFF; assign b = 64'h01DFFFFFFFFFFFFF;

    #10 $display("\n2**-80 * 2**-995:");
    #10 assign a = 64'h3AF0000000000000; assign b = 64'h01C0000000000000;
    #10 assign a = 64'h3AFFFFFFFFFFFFFF; assign b = 64'h01CFFFFFFFFFFFFF;

    #10 $display("\n2**-79 * 2**-996:");
    #10 assign a = 64'h3B00000000000000; assign b = 64'h01B0000000000000;
    #10 assign a = 64'h3B0FFFFFFFFFFFFF; assign b = 64'h01BFFFFFFFFFFFFF;

    #10 $display("\n2**-78 * 2**-997:");
    #10 assign a = 64'h3B10000000000000; assign b = 64'h01A0000000000000;
    #10 assign a = 64'h3B1FFFFFFFFFFFFF; assign b = 64'h01AFFFFFFFFFFFFF;

    #10 $display("\n2**-77 * 2**-998:");
    #10 assign a = 64'h3B20000000000000; assign b = 64'h0190000000000000;
    #10 assign a = 64'h3B2FFFFFFFFFFFFF; assign b = 64'h019FFFFFFFFFFFFF;

    #10 $display("\n2**-76 * 2**-999:");
    #10 assign a = 64'h3B30000000000000; assign b = 64'h0180000000000000;
    #10 assign a = 64'h3B3FFFFFFFFFFFFF; assign b = 64'h018FFFFFFFFFFFFF;

    #10 $display("\n2**-75 * 2**-1000:");
    #10 assign a = 64'h3B40000000000000; assign b = 64'h0170000000000000;
    #10 assign a = 64'h3B4FFFFFFFFFFFFF; assign b = 64'h017FFFFFFFFFFFFF;

    #10 $display("\n2**-74 * 2**-1001:");
    #10 assign a = 64'h3B50000000000000; assign b = 64'h0160000000000000;
    #10 assign a = 64'h3B5FFFFFFFFFFFFF; assign b = 64'h016FFFFFFFFFFFFF;

    #10 $display("\n2**-73 * 2**-1002:");
    #10 assign a = 64'h3B60000000000000; assign b = 64'h0150000000000000;
    #10 assign a = 64'h3B6FFFFFFFFFFFFF; assign b = 64'h015FFFFFFFFFFFFF;

    #10 $display("\n2**-72 * 2**-1003:");
    #10 assign a = 64'h3B70000000000000; assign b = 64'h0140000000000000;
    #10 assign a = 64'h3B7FFFFFFFFFFFFF; assign b = 64'h014FFFFFFFFFFFFF;

    #10 $display("\n2**-71 * 2**-1004:");
    #10 assign a = 64'h3B80000000000000; assign b = 64'h0130000000000000;
    #10 assign a = 64'h3B8FFFFFFFFFFFFF; assign b = 64'h013FFFFFFFFFFFFF;

    #10 $display("\n2**-70 * 2**-1005:");
    #10 assign a = 64'h3B90000000000000; assign b = 64'h0120000000000000;
    #10 assign a = 64'h3B9FFFFFFFFFFFFF; assign b = 64'h012FFFFFFFFFFFFF;

    #10 $display("\n2**-69 * 2**-1006:");
    #10 assign a = 64'h3BA0000000000000; assign b = 64'h0110000000000000;
    #10 assign a = 64'h3BAFFFFFFFFFFFFF; assign b = 64'h011FFFFFFFFFFFFF;

    #10 $display("\n2**-68 * 2**-1007:");
    #10 assign a = 64'h3BB0000000000000; assign b = 64'h0100000000000000;
    #10 assign a = 64'h3BBFFFFFFFFFFFFF; assign b = 64'h010FFFFFFFFFFFFF;

    #10 $display("\n2**-67 * 2**-1008:");
    #10 assign a = 64'h3BC0000000000000; assign b = 64'h00F0000000000000;
    #10 assign a = 64'h3BCFFFFFFFFFFFFF; assign b = 64'h00FFFFFFFFFFFFFF;

    #10 $display("\n2**-66 * 2**-1009:");
    #10 assign a = 64'h3BD0000000000000; assign b = 64'h00E0000000000000;
    #10 assign a = 64'h3BDFFFFFFFFFFFFF; assign b = 64'h00EFFFFFFFFFFFFF;

    #10 $display("\n2**-65 * 2**-1010:");
    #10 assign a = 64'h3BE0000000000000; assign b = 64'h00D0000000000000;
    #10 assign a = 64'h3BEFFFFFFFFFFFFF; assign b = 64'h00DFFFFFFFFFFFFF;

    #10 $display("\n2**-64 * 2**-1011:");
    #10 assign a = 64'h3BF0000000000000; assign b = 64'h00C0000000000000;
    #10 assign a = 64'h3BFFFFFFFFFFFFFF; assign b = 64'h00CFFFFFFFFFFFFF;

    #10 $display("\n2**-63 * 2**-1012:");
    #10 assign a = 64'h3C00000000000000; assign b = 64'h00B0000000000000;
    #10 assign a = 64'h3C0FFFFFFFFFFFFF; assign b = 64'h00BFFFFFFFFFFFFF;

    #10 $display("\n2**-62 * 2**-1013:");
    #10 assign a = 64'h3C10000000000000; assign b = 64'h00A0000000000000;
    #10 assign a = 64'h3C1FFFFFFFFFFFFF; assign b = 64'h00AFFFFFFFFFFFFF;

    #10 $display("\n2**-61 * 2**-1014:");
    #10 assign a = 64'h3C20000000000000; assign b = 64'h0090000000000000;
    #10 assign a = 64'h3C2FFFFFFFFFFFFF; assign b = 64'h009FFFFFFFFFFFFF;

    #10 $display("\n2**-60 * 2**-1015:");
    #10 assign a = 64'h3C30000000000000; assign b = 64'h0080000000000000;
    #10 assign a = 64'h3C3FFFFFFFFFFFFF; assign b = 64'h008FFFFFFFFFFFFF;

    #10 $display("\n2**-59 * 2**-1016:");
    #10 assign a = 64'h3C40000000000000; assign b = 64'h0070000000000000;
    #10 assign a = 64'h3C4FFFFFFFFFFFFF; assign b = 64'h007FFFFFFFFFFFFF;

    #10 $display("\n2**-58 * 2**-1017:");
    #10 assign a = 64'h3C50000000000000; assign b = 64'h0060000000000000;
    #10 assign a = 64'h3C5FFFFFFFFFFFFF; assign b = 64'h006FFFFFFFFFFFFF;

    #10 $display("\n2**-57 * 2**-1018:");
    #10 assign a = 64'h3C60000000000000; assign b = 64'h0050000000000000;
    #10 assign a = 64'h3C6FFFFFFFFFFFFF; assign b = 64'h005FFFFFFFFFFFFF;

    #10 $display("\n2**-56 * 2**-1019:");
    #10 assign a = 64'h3C70000000000000; assign b = 64'h0040000000000000;
    #10 assign a = 64'h3C7FFFFFFFFFFFFF; assign b = 64'h004FFFFFFFFFFFFF;

    #10 $display("\n2**-55 * 2**-1020:");
    #10 assign a = 64'h3C80000000000000; assign b = 64'h0030000000000000;
    #10 assign a = 64'h3C8FFFFFFFFFFFFF; assign b = 64'h003FFFFFFFFFFFFF;

    #10 $display("\n2**-54 * 2**-1021:");
    #10 assign a = 64'h3C90000000000000; assign b = 64'h0020000000000000;
    #10 assign a = 64'h3C9FFFFFFFFFFFFF; assign b = 64'h002FFFFFFFFFFFFF;

    #10 $display("\n2**-53 * 2**-1022:");
    #10 assign a = 64'h3CA0000000000000; assign b = 64'h0010000000000000;
    #10 assign a = 64'h3CAFFFFFFFFFFFFF; assign b = 64'h001FFFFFFFFFFFFF;

    #10 $display("\n2**-52 * 2**-1023:");
    #10 assign a = 64'h3CB0000000000000; assign b = 64'h0008000000000000;
    #10 assign a = 64'h3CBFFFFFFFFFFFFF; assign b = 64'h000FFFFFFFFFFFFF;

    #10 $display("\n2**-51 * 2**-1024:");
    #10 assign a = 64'h3CC0000000000000; assign b = 64'h0004000000000000;
    #10 assign a = 64'h3CCFFFFFFFFFFFFF; assign b = 64'h0007FFFFFFFFFFFF;

    #10 $display("\n2**-50 * 2**-1025:");
    #10 assign a = 64'h3CD0000000000000; assign b = 64'h0002000000000000;
    #10 assign a = 64'h3CDFFFFFFFFFFFFF; assign b = 64'h0003FFFFFFFFFFFF;

    #10 $display("\n2**-49 * 2**-1026:");
    #10 assign a = 64'h3CE0000000000000; assign b = 64'h0001000000000000;
    #10 assign a = 64'h3CEFFFFFFFFFFFFF; assign b = 64'h0001FFFFFFFFFFFF;

    #10 $display("\n2**-48 * 2**-1027:");
    #10 assign a = 64'h3CF0000000000000; assign b = 64'h0000800000000000;
    #10 assign a = 64'h3CFFFFFFFFFFFFFF; assign b = 64'h0000FFFFFFFFFFFF;

    #10 $display("\n2**-47 * 2**-1028:");
    #10 assign a = 64'h3D00000000000000; assign b = 64'h0000400000000000;
    #10 assign a = 64'h3D0FFFFFFFFFFFFF; assign b = 64'h00007FFFFFFFFFFF;

    #10 $display("\n2**-46 * 2**-1029:");
    #10 assign a = 64'h3D10000000000000; assign b = 64'h0000200000000000;
    #10 assign a = 64'h3D1FFFFFFFFFFFFF; assign b = 64'h00003FFFFFFFFFFF;

    #10 $display("\n2**-45 * 2**-1030:");
    #10 assign a = 64'h3D20000000000000; assign b = 64'h0000100000000000;
    #10 assign a = 64'h3D2FFFFFFFFFFFFF; assign b = 64'h00001FFFFFFFFFFF;

    #10 $display("\n2**-44 * 2**-1031:");
    #10 assign a = 64'h3D30000000000000; assign b = 64'h0000080000000000;
    #10 assign a = 64'h3D3FFFFFFFFFFFFF; assign b = 64'h00000FFFFFFFFFFF;

    #10 $display("\n2**-43 * 2**-1032:");
    #10 assign a = 64'h3D40000000000000; assign b = 64'h0000040000000000;
    #10 assign a = 64'h3D4FFFFFFFFFFFFF; assign b = 64'h000007FFFFFFFFFF;

    #10 $display("\n2**-42 * 2**-1033:");
    #10 assign a = 64'h3D50000000000000; assign b = 64'h0000020000000000;
    #10 assign a = 64'h3D5FFFFFFFFFFFFF; assign b = 64'h000003FFFFFFFFFF;

    #10 $display("\n2**-41 * 2**-1034:");
    #10 assign a = 64'h3D60000000000000; assign b = 64'h0000010000000000;
    #10 assign a = 64'h3D6FFFFFFFFFFFFF; assign b = 64'h000001FFFFFFFFFF;

    #10 $display("\n2**-40 * 2**-1035:");
    #10 assign a = 64'h3D70000000000000; assign b = 64'h0000008000000000;
    #10 assign a = 64'h3D7FFFFFFFFFFFFF; assign b = 64'h000000FFFFFFFFFF;

    #10 $display("\n2**-39 * 2**-1036:");
    #10 assign a = 64'h3D80000000000000; assign b = 64'h0000004000000000;
    #10 assign a = 64'h3D8FFFFFFFFFFFFF; assign b = 64'h0000007FFFFFFFFF;

    #10 $display("\n2**-38 * 2**-1037:");
    #10 assign a = 64'h3D90000000000000; assign b = 64'h0000002000000000;
    #10 assign a = 64'h3D9FFFFFFFFFFFFF; assign b = 64'h0000003FFFFFFFFF;

    #10 $display("\n2**-37 * 2**-1038:");
    #10 assign a = 64'h3DA0000000000000; assign b = 64'h0000001000000000;
    #10 assign a = 64'h3DAFFFFFFFFFFFFF; assign b = 64'h0000001FFFFFFFFF;

    #10 $display("\n2**-36 * 2**-1039:");
    #10 assign a = 64'h3DB0000000000000; assign b = 64'h0000000800000000;
    #10 assign a = 64'h3DBFFFFFFFFFFFFF; assign b = 64'h0000000FFFFFFFFF;

    #10 $display("\n2**-35 * 2**-1040:");
    #10 assign a = 64'h3DC0000000000000; assign b = 64'h0000000400000000;
    #10 assign a = 64'h3DCFFFFFFFFFFFFF; assign b = 64'h00000007FFFFFFFF;

    #10 $display("\n2**-34 * 2**-1041:");
    #10 assign a = 64'h3DD0000000000000; assign b = 64'h0000000200000000;
    #10 assign a = 64'h3DDFFFFFFFFFFFFF; assign b = 64'h00000003FFFFFFFF;

    #10 $display("\n2**-33 * 2**-1042:");
    #10 assign a = 64'h3DE0000000000000; assign b = 64'h0000000100000000;
    #10 assign a = 64'h3DEFFFFFFFFFFFFF; assign b = 64'h00000001FFFFFFFF;

    #10 $display("\n2**-32 * 2**-1043:");
    #10 assign a = 64'h3DF0000000000000; assign b = 64'h0000000080000000;
    #10 assign a = 64'h3DFFFFFFFFFFFFFF; assign b = 64'h00000000FFFFFFFF;

    #10 $display("\n2**-31 * 2**-1044:");
    #10 assign a = 64'h3E00000000000000; assign b = 64'h0000000040000000;
    #10 assign a = 64'h3E0FFFFFFFFFFFFF; assign b = 64'h000000007FFFFFFF;

    #10 $display("\n2**-30 * 2**-1045:");
    #10 assign a = 64'h3E10000000000000; assign b = 64'h0000000020000000;
    #10 assign a = 64'h3E1FFFFFFFFFFFFF; assign b = 64'h000000003FFFFFFF;

    #10 $display("\n2**-29 * 2**-1046:");
    #10 assign a = 64'h3E20000000000000; assign b = 64'h0000000010000000;
    #10 assign a = 64'h3E2FFFFFFFFFFFFF; assign b = 64'h000000001FFFFFFF;

    #10 $display("\n2**-28 * 2**-1047:");
    #10 assign a = 64'h3E30000000000000; assign b = 64'h0000000008000000;
    #10 assign a = 64'h3E3FFFFFFFFFFFFF; assign b = 64'h000000000FFFFFFF;

    #10 $display("\n2**-27 * 2**-1048:");
    #10 assign a = 64'h3E40000000000000; assign b = 64'h0000000004000000;
    #10 assign a = 64'h3E4FFFFFFFFFFFFF; assign b = 64'h0000000007FFFFFF;

    #10 $display("\n2**-26 * 2**-1049:");
    #10 assign a = 64'h3E50000000000000; assign b = 64'h0000000002000000;
    #10 assign a = 64'h3E5FFFFFFFFFFFFF; assign b = 64'h0000000003FFFFFF;

    #10 $display("\n2**-25 * 2**-1050:");
    #10 assign a = 64'h3E60000000000000; assign b = 64'h0000000001000000;
    #10 assign a = 64'h3E6FFFFFFFFFFFFF; assign b = 64'h0000000001FFFFFF;

    #10 $display("\n2**-24 * 2**-1051:");
    #10 assign a = 64'h3E70000000000000; assign b = 64'h0000000000800000;
    #10 assign a = 64'h3E7FFFFFFFFFFFFF; assign b = 64'h0000000000FFFFFF;

    #10 $display("\n2**-23 * 2**-1052:");
    #10 assign a = 64'h3E80000000000000; assign b = 64'h0000000000400000;
    #10 assign a = 64'h3E8FFFFFFFFFFFFF; assign b = 64'h00000000007FFFFF;

    #10 $display("\n2**-22 * 2**-1053:");
    #10 assign a = 64'h3E90000000000000; assign b = 64'h0000000000200000;
    #10 assign a = 64'h3E9FFFFFFFFFFFFF; assign b = 64'h00000000003FFFFF;

    #10 $display("\n2**-21 * 2**-1054:");
    #10 assign a = 64'h3EA0000000000000; assign b = 64'h0000000000100000;
    #10 assign a = 64'h3EAFFFFFFFFFFFFF; assign b = 64'h00000000001FFFFF;

    #10 $display("\n2**-20 * 2**-1055:");
    #10 assign a = 64'h3EB0000000000000; assign b = 64'h0000000000080000;
    #10 assign a = 64'h3EBFFFFFFFFFFFFF; assign b = 64'h00000000000FFFFF;

    #10 $display("\n2**-19 * 2**-1056:");
    #10 assign a = 64'h3EC0000000000000; assign b = 64'h0000000000040000;
    #10 assign a = 64'h3ECFFFFFFFFFFFFF; assign b = 64'h000000000007FFFF;

    #10 $display("\n2**-18 * 2**-1057:");
    #10 assign a = 64'h3ED0000000000000; assign b = 64'h0000000000020000;
    #10 assign a = 64'h3EDFFFFFFFFFFFFF; assign b = 64'h000000000003FFFF;

    #10 $display("\n2**-17 * 2**-1058:");
    #10 assign a = 64'h3EE0000000000000; assign b = 64'h0000000000010000;
    #10 assign a = 64'h3EEFFFFFFFFFFFFF; assign b = 64'h000000000001FFFF;

    #10 $display("\n2**-16 * 2**-1059:");
    #10 assign a = 64'h3EF0000000000000; assign b = 64'h0000000000008000;
    #10 assign a = 64'h3EFFFFFFFFFFFFFF; assign b = 64'h000000000000FFFF;

    #10 $display("\n2**-15 * 2**-1060:");
    #10 assign a = 64'h3F00000000000000; assign b = 64'h0000000000004000;
    #10 assign a = 64'h3F0FFFFFFFFFFFFF; assign b = 64'h0000000000007FFF;

    #10 $display("\n2**-14 * 2**-1061:");
    #10 assign a = 64'h3F10000000000000; assign b = 64'h0000000000002000;
    #10 assign a = 64'h3F1FFFFFFFFFFFFF; assign b = 64'h0000000000003FFF;

    #10 $display("\n2**-13 * 2**-1062:");
    #10 assign a = 64'h3F20000000000000; assign b = 64'h0000000000001000;
    #10 assign a = 64'h3F2FFFFFFFFFFFFF; assign b = 64'h0000000000001FFF;

    #10 $display("\n2**-12 * 2**-1063:");
    #10 assign a = 64'h3F30000000000000; assign b = 64'h0000000000000800;
    #10 assign a = 64'h3F3FFFFFFFFFFFFF; assign b = 64'h0000000000000FFF;

    #10 $display("\n2**-11 * 2**-1064:");
    #10 assign a = 64'h3F40000000000000; assign b = 64'h0000000000000400;
    #10 assign a = 64'h3F4FFFFFFFFFFFFF; assign b = 64'h00000000000007FF;

    #10 $display("\n2**-10 * 2**-1065:");
    #10 assign a = 64'h3F50000000000000; assign b = 64'h0000000000000200;
    #10 assign a = 64'h3F5FFFFFFFFFFFFF; assign b = 64'h00000000000003FF;

    #10 $display("\n2**-9 * 2**-1066:");
    #10 assign a = 64'h3F60000000000000; assign b = 64'h0000000000000100;
    #10 assign a = 64'h3F6FFFFFFFFFFFFF; assign b = 64'h00000000000001FF;

    #10 $display("\n2**-8 * 2**-1067:");
    #10 assign a = 64'h3F70000000000000; assign b = 64'h0000000000000080;
    #10 assign a = 64'h3F7FFFFFFFFFFFFF; assign b = 64'h00000000000000FF;

    #10 $display("\n2**-7 * 2**-1068:");
    #10 assign a = 64'h3F80000000000000; assign b = 64'h0000000000000040;
    #10 assign a = 64'h3F8FFFFFFFFFFFFF; assign b = 64'h000000000000007F;

    #10 $display("\n2**-6 * 2**-1069:");
    #10 assign a = 64'h3F90000000000000; assign b = 64'h0000000000000020;
    #10 assign a = 64'h3F9FFFFFFFFFFFFF; assign b = 64'h000000000000003F;

    #10 $display("\n2**-5 * 2**-1070:");
    #10 assign a = 64'h3FA0000000000000; assign b = 64'h0000000000000010;
    #10 assign a = 64'h3FAFFFFFFFFFFFFF; assign b = 64'h000000000000001F;

    #10 $display("\n2**-4 * 2**-1071:");
    #10 assign a = 64'h3FB0000000000000; assign b = 64'h0000000000000008;
    #10 assign a = 64'h3FBFFFFFFFFFFFFF; assign b = 64'h000000000000000F;

    #10 $display("\n2**-3 * 2**-1072:");
    #10 assign a = 64'h3FC0000000000000; assign b = 64'h0000000000000004;
    #10 assign a = 64'h3FCFFFFFFFFFFFFF; assign b = 64'h0000000000000007;

    #10 $display("\n2**-2 * 2**-1073:");
    #10 assign a = 64'h3FD0000000000000; assign b = 64'h0000000000000002;
    #10 assign a = 64'h3FDFFFFFFFFFFFFF; assign b = 64'h0000000000000003;

    #10 $display("\n2**-1 * 2**-1074:");
    #10 assign a = 64'h3FE0000000000000; assign b = 64'h0000000000000001;
    #10 assign a = 64'h3FEFFFFFFFFFFFFF; assign b = 64'h0000000000000001;

//    #10 $display("\n20 * 20:"); // 1.0100000000 * 2**4 or 0x4D00
//    #10 assign a = 16'h4D00; assign b = 16'h4D00; // 1.1001000000 x 2**8 or 0x5E40
//
//    #10 $display("\n400 * PI:"); // PI = 1.1001001000 * 2**1
//    #10 assign a = 16'h5E40; assign b = 16'h4248; // 1.0011101000 * 2**10 or 0x64E8

    #20 $display("\nEnd of tests : %t", $time);
    #20 $stop;
  end

  fp_mul #(NEXP, NSIG) inst1(
  .a(a),
  .b(b),
  .p(p),
  .pFlags(flags)
  );
endmodule
